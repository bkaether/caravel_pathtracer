
//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v5.v 
module mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features; 
//       please enable Verilog2001 in the flow!

module mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers
   
    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC
   
    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_genreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_genreg_v1 (clk, en, arst, srst, d, z);
    parameter integer width   = 1;
    parameter integer ph_clk  = 1;
    parameter integer ph_en   = 1;
    parameter integer ph_arst = 0;
    parameter integer ph_srst = 1;
    parameter         has_en  = 1'b1;

    input clk;
    input en;
    input arst;
    input srst;
    input      [width-1:0] d;
    output reg [width-1:0] z;

    //  Generate parameters
    //  ph_clk | ph_arst | has_en     Label:
    //    1        1          1       GEN_CLK1_ARST1_EN1
    //    1        1          0       GEN_CLK1_ARST1_EN0
    //    1        0          1       GEN_CLK1_ARST0_EN1
    //    1        0          0       GEN_CLK1_ARST0_EN0
    //    0        1          1       GEN_CLK0_ARST1_EN1
    //    0        1          0       GEN_CLK0_ARST1_EN0
    //    0        0          1       GEN_CLK0_ARST0_EN1
    //    0        0          0       GEN_CLK0_ARST0_EN0
    
    generate 
      // Pos edge clock, pos edge async reset, has enable
      if (ph_clk == 1 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK1_ARST1_EN1
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST1_EN1

      // Pos edge clock, pos edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK1_ARST1_EN0
        always @(posedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST1_EN0

      // Pos edge clock, neg edge async reset, has enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK1_ARST0_EN1
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK1_ARST0_EN1

      // Pos edge clock, neg edge async reset, no enable
      else if (ph_clk == 1 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK1_ARST0_EN0
        always @(posedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK1_ARST0_EN0


      // Neg edge clock, pos edge async reset, has enable
      if (ph_clk == 0 & ph_arst == 1 & has_en == 1)
      begin: GEN_CLK0_ARST1_EN1
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST1_EN1

      // Neg edge clock, pos edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 1 & has_en == 0)
      begin: GEN_CLK0_ARST1_EN0
        always @(negedge clk or posedge arst)
          if (arst == 1'b1)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST1_EN0

      // Neg edge clock, neg edge async reset, has enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 1)
      begin: GEN_CLK0_ARST0_EN1
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else if (en == $unsigned(ph_en))
            z <= d;
      end  //GEN_CLK0_ARST0_EN1

      // Neg edge clock, neg edge async reset, no enable
      else if (ph_clk == 0 & ph_arst == 0 & has_en == 0)
      begin: GEN_CLK0_ARST0_EN0
        always @(negedge clk or negedge arst)
          if (arst == 1'b0)
            z <= {width{1'b0}};
          else if (srst == $unsigned(ph_srst))
            z <= {width{1'b0}};
          else
            z <= d;
      end  //GEN_CLK0_ARST0_EN0
    endgenerate
endmodule


//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_fifo_wait_core_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

/*
 *            _________________________________________________
 * WRITER    |                                                 |   READER
 *           |               ccs_fifo_wait_core                |
 *           |             _____________________               |
 *        --<|  din_rdy --<|  ---------------- <|--- dout_rdy <|---
 *           |             |       FIFO         |              |
 *        ---|> din_vld ---|> ----------------  |>-- dout_vld  |>--
 *        ---|>     din ---|> ----------------  |>-- dout      |>--
 *           |             |____________________|              |
 *           |_________________________________________________|
 *
 *    rdy    - can be considered as a notFULL signal
 *    vld    - can be considered as a notEMPTY signal
 *    is_idle - clk can be safely gated
 *
 * Change History:
 *    2019-01-24 - Add assertion to verify rdy signal behavior under reset.
 *                 Fix bug in that behavior.
 */

module ccs_fifo_wait_core_v5 (clk, en, arst, srst, din_vld, din_rdy, din, dout_vld, dout_rdy, dout, sd, is_idle);

    parameter integer rscid    = 0;     // resource ID
    parameter integer width    = 8;     // fifo width
    parameter integer sz_width = 8;     // size of port for elements in fifo
    parameter integer fifo_sz  = 8;     // fifo depth
    parameter integer ph_clk   = 1;  // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1;  // clock enable polarity
    parameter integer ph_arst  = 1;  // async reset polarity
    parameter integer ph_srst  = 1;  // sync reset polarity
    parameter integer ph_log2  = 3;     // log2(fifo_sz)

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 din_vld;    // writer has valid data 
    output                din_rdy;    // fifo ready for data (not full)
    input  [width-1:0]    din;
    output                dout_vld;   // fifo has valid data (not empty)
    input                 dout_rdy;   // reader ready for data
    output [width-1:0]    dout;
    output [sz_width-1:0] sd; 
    output                is_idle;

    localparam integer fifo_b  = width * fifo_sz;
    localparam integer fifo_mx = (fifo_sz > 0) ? (fifo_sz-1) : 0 ;
    localparam integer fifo_mx_over_8 = fifo_mx / 8 ;

    reg      [fifo_mx:0] stat_pre;
    wire     [fifo_mx:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [fifo_mx:0] en_l;
    reg      [fifo_mx_over_8:0] en_l_s;

    reg      [width-1:0] buff_nxt;

    reg                  stat_nxt;
    reg                  stat_behind;
    reg                  stat_ahead;
    reg                  en_l_var;

    integer              i;
    genvar               eni;

    wire [32:0]          size_t;
    reg  [31:0]          count;
    reg  [31:0]          count_t;
    reg  [32:0]          n_elem;
    // synopsys translate_off
    reg  [31:0]          peak;
    initial
    begin
      count = 32'b0;
      peak  = 32'b0;
    end
    // synopsys translate_on
  wire din_rdy_drv  ;
  wire dout_vld_drv ;
    wire                 active;
    wire                 din_vld_int;
    wire                 hs_init;

    //assign din_rdy  = din_rdy_drv;    // dout_rdy | (~stat[0] & hs_init);   // original
    assign din_rdy = (fifo_sz > 0) ? (~stat[0] | dout_rdy) && hs_init : dout_rdy ;       // experiment
 
    assign dout_vld = dout_vld_drv;
    assign is_idle = (~((din_vld && din_rdy) || (dout_vld && dout_rdy))) && hs_init;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
    assign din_vld_int = din_vld & hs_init;
    // KH assign active = din_vld_int | dout_rdy; // (din_vld & ~din_rdy) | (dout_rdy & ~dout_vld);
    assign active =   (din_vld_int & din_rdy_drv) | (dout_rdy & dout_vld_drv);

      assign din_rdy_drv = dout_rdy | (~stat[0] & hs_init);
      assign dout_vld_drv = din_vld_int | stat[fifo_sz-1];

      assign size_t = (count - {31'b0 , (dout_rdy & stat[fifo_sz-1])}) + { 31'b0, din_vld_int};
      assign sd = size_t[sz_width-1:0];

      assign dout = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : din;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          stat_behind = (i != 0) ? stat[i-1] : 1'b0;
          stat_ahead  = (i != (fifo_sz-1)) ? stat[i+1] : 1'b1;

          // Determine if this buffer element will have data
          stat_nxt = stat_ahead &                       // valid element ahead of this one (or head)
                       (stat_behind                     // valid element behind this one
                         | (stat[i] & (~dout_rdy))      // valid element and output not ready (in use, no tx)
                         | (stat[i] & din_vld_int)      // valid element and input has data
                         | (din_vld_int  & (~dout_rdy)) // input has data and output not ready
                       );
          stat_pre[i] = stat_nxt;

          if (dout_rdy & stat_behind )
          begin
            // pop n shift
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
            en_l_var = 1'b1;
          end
          else if (din_vld_int & stat_nxt & ~((~dout_rdy) & stat[i]))
          begin
            // update tail with input data
            buff_nxt = din;
            en_l_var = 1'b1;
          end
          else
          begin
            // no-op, disable register
            buff_nxt = din; // Don't care input to disabled flop
            en_l_var = 1'b0;
          end
          buff_pre[width*i+:width] = buff_nxt[0+:width];
             
          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          if ((stat_ahead == 1'b1) & (stat[i] == 1'b0)) 
            //found tail, update the number of elements for count
            n_elem = ($unsigned(fifo_sz) - 1) - $unsigned(i);
        end //for loop

        // Enable for stat registers (partitioned into banks of eight)
        // Take care of the head first
        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en & active;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = en | ~active;

        // Now every eight
        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if (($unsigned(i)%8) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]) & (active);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]) | ~(active);
          end
        end
        
        // Update count and peak
        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = fifo_sz;
        else 
          count_t = n_elem[31:0];
        count = count_t;
        // synopsys translate_off
        if ( peak < count )
          peak = count;
        // synopsys translate_on
      end //FIFOPROC

      // Handshake valid after reset
      ccs_genreg_v1
      #(
        .width   (1),
        .ph_clk  (ph_clk),
        .ph_en   (1),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .has_en  (1'b0)
      )
      HS_INIT_REG
      (
        .clk     (clk),
        .en      (1'b1),
        .arst    (arst),
        .srst    (srst),
        .d       (1'b1),
        .z       (hs_init)
      );

      // Buffer and status registers
      for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
      begin: GEN_REGS
        ccs_genreg_v1
        #(
          .width   (1),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        STATREG
        (
          .clk     (clk),
          .en      (en_l_s[eni/8]),
          .arst    (arst),
          .srst    (srst),
          .d       (stat_pre[eni]),
          .z       (stat[eni])
        );

        ccs_genreg_v1
        #(
          .width   (width),
          .ph_clk  (ph_clk),
          .ph_en   (ph_en),
          .ph_arst (ph_arst),
          .ph_srst (ph_srst),
          .has_en  (1'b1)
        )
        BUFREG
        (
          .clk     (clk),
          .en      (en_l[eni]),
          .arst    (arst),
          .srst    (srst),
          .d       (buff_pre[width*eni+:width]),
          .z       (buff[width*eni+:width])
        );
      end

    end
    else
    begin: FEED_THRU
      assign din_rdy_drv  = dout_rdy;
      assign dout_vld_drv = din_vld;
      assign dout     = din;
      // non-blocking is not II=1 when fifo_sz=0
      assign sd = {{(sz_width-1){1'b0}}, (din_vld & ~dout_rdy)};
    end
    endgenerate

`ifdef RDY_ASRT 
    generate
    if (ph_clk==1) 
    begin: POS_CLK_ASSERT

       property rdyAsrt ;
         @(posedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Pos: assert property(rdyAsrt);

    end else if (ph_clk==0) 
    begin: NEG_CLK_ASSERT

       property rdyAsrt ;
         @(negedge clk) ((srst==ph_srst) || (arst==ph_arst)) |=> (din_rdy==0);
       endproperty
       a1Neg: assert property(rdyAsrt);

    end
    endgenerate

`endif
   
endmodule



//------> /cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_pipe_v5.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
/*
 *
 *            _______________________________________________
 * WRITER    |                                              |          READER
 *           |                 ccs_pipe                     |
 *           |            ______________________            |
 *        --<| din_rdy --<|  ---------------- <|---dout_rdy<|---
 *           |            |       FIFO         |            |
 *        ---|>din_vld ---|> ----------------  |>--dout_vld |>--
 *        ---|>din -------|> ----------------  |> -----dout |>--
 *           |            |____________________|            |
 *           |______________________________________________|
 *
 *    din_rdy     - can be considered as a notFULL signal
 *    dout_vld    - can be considered as a notEMPTY signal
 *    write_stall - an internal debug signal formed from din_vld & !din_rdy
 *    read_stall  - an internal debug signal formed from dout_rdy & !dout_vld
 *    is_idle     - indicates the clock can be safely gated
 */

module ccs_pipe_v5 (clk, en, arst, srst, din_rdy, din_vld, din, dout_rdy, dout_vld, dout, sz, sz_req, is_idle);

    parameter integer rscid    = 0; // resource ID
    parameter integer width    = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz  = 8; // fifo depth
    parameter integer log2_sz  = 3; // log2(fifo_sz)
    parameter integer ph_clk   = 1; // clock polarity 1=rising edge, 0=falling edge
    parameter integer ph_en    = 1; // clock enable polarity
    parameter integer ph_arst  = 1; // async reset polarity
    parameter integer ph_srst  = 1; // sync reset polarity

    // clock 
    input              clk;
    input              en;
    input              arst;
    input              srst;

    // writer
    output             din_rdy;
    input              din_vld;
    input  [width-1:0] din;

    // reader
    input              dout_rdy;
    output             dout_vld;
    output [width-1:0] dout;

    // size
    output [sz_width-1:0] sz;
    input                 sz_req;
    output                is_idle;
   
    // synopsys translate_off
    wire   write_stall;
    wire   read_stall;
    assign write_stall = din_vld & !din_rdy;
    assign read_stall  = dout_rdy & !dout_vld;
    // synopsys translate_on

    ccs_fifo_wait_core_v5
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz)
    )
    FIFO
    (
        .clk      (clk),
        .en       (en),
        .arst     (arst),
        .srst     (srst),
        .din_vld  (din_vld),
        .din_rdy  (din_rdy),
        .din      (din),
        .dout_vld (dout_vld),
        .dout_rdy (dout_rdy),
        .dout     (dout),
        .sd       (sz),
        .is_idle  (is_idle)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   bkaether@iron-02
//  Generated date: Sun Jun  2 15:17:10 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ParamsDeserializer_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, for_C_41_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input for_C_41_tr0;


  // FSM State Type Declaration for ParamsDeserializer_run_run_fsm_1
  parameter
    run_rlp_C_0 = 7'd0,
    main_C_0 = 7'd1,
    main_C_1 = 7'd2,
    main_C_2 = 7'd3,
    main_C_3 = 7'd4,
    main_C_4 = 7'd5,
    main_C_5 = 7'd6,
    main_C_6 = 7'd7,
    main_C_7 = 7'd8,
    main_C_8 = 7'd9,
    main_C_9 = 7'd10,
    main_C_10 = 7'd11,
    main_C_11 = 7'd12,
    main_C_12 = 7'd13,
    main_C_13 = 7'd14,
    main_C_14 = 7'd15,
    main_C_15 = 7'd16,
    main_C_16 = 7'd17,
    main_C_17 = 7'd18,
    main_C_18 = 7'd19,
    main_C_19 = 7'd20,
    main_C_20 = 7'd21,
    main_C_21 = 7'd22,
    main_C_22 = 7'd23,
    main_C_23 = 7'd24,
    main_C_24 = 7'd25,
    main_C_25 = 7'd26,
    main_C_26 = 7'd27,
    main_C_27 = 7'd28,
    main_C_28 = 7'd29,
    main_C_29 = 7'd30,
    main_C_30 = 7'd31,
    main_C_31 = 7'd32,
    main_C_32 = 7'd33,
    main_C_33 = 7'd34,
    main_C_34 = 7'd35,
    main_C_35 = 7'd36,
    main_C_36 = 7'd37,
    main_C_37 = 7'd38,
    main_C_38 = 7'd39,
    main_C_39 = 7'd40,
    main_C_40 = 7'd41,
    main_C_41 = 7'd42,
    main_C_42 = 7'd43,
    main_C_43 = 7'd44,
    main_C_44 = 7'd45,
    main_C_45 = 7'd46,
    for_C_0 = 7'd47,
    for_C_1 = 7'd48,
    for_C_2 = 7'd49,
    for_C_3 = 7'd50,
    for_C_4 = 7'd51,
    for_C_5 = 7'd52,
    for_C_6 = 7'd53,
    for_C_7 = 7'd54,
    for_C_8 = 7'd55,
    for_C_9 = 7'd56,
    for_C_10 = 7'd57,
    for_C_11 = 7'd58,
    for_C_12 = 7'd59,
    for_C_13 = 7'd60,
    for_C_14 = 7'd61,
    for_C_15 = 7'd62,
    for_C_16 = 7'd63,
    for_C_17 = 7'd64,
    for_C_18 = 7'd65,
    for_C_19 = 7'd66,
    for_C_20 = 7'd67,
    for_C_21 = 7'd68,
    for_C_22 = 7'd69,
    for_C_23 = 7'd70,
    for_C_24 = 7'd71,
    for_C_25 = 7'd72,
    for_C_26 = 7'd73,
    for_C_27 = 7'd74,
    for_C_28 = 7'd75,
    for_C_29 = 7'd76,
    for_C_30 = 7'd77,
    for_C_31 = 7'd78,
    for_C_32 = 7'd79,
    for_C_33 = 7'd80,
    for_C_34 = 7'd81,
    for_C_35 = 7'd82,
    for_C_36 = 7'd83,
    for_C_37 = 7'd84,
    for_C_38 = 7'd85,
    for_C_39 = 7'd86,
    for_C_40 = 7'd87,
    for_C_41 = 7'd88;

  reg [6:0] state_var;
  reg [6:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ParamsDeserializer_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 7'b0000010;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b0000011;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b0000100;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 7'b0000101;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 7'b0000110;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 7'b0000111;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 7'b0001000;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 7'b0001001;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 7'b0001010;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 7'b0001011;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 7'b0001100;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 7'b0001101;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 7'b0001110;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 7'b0001111;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 7'b0010000;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 7'b0010001;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 7'b0010010;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 7'b0010011;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 7'b0010100;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 7'b0010101;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 7'b0010110;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 7'b0010111;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 7'b0011000;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 7'b0011001;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 7'b0011010;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 7'b0011011;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 7'b0011100;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 7'b0011101;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 7'b0011110;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 7'b0011111;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 7'b0100000;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 7'b0100001;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 7'b0100010;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 7'b0100011;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 7'b0100100;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 7'b0100101;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 7'b0100110;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 7'b0100111;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 7'b0101000;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 7'b0101001;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 7'b0101010;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 7'b0101011;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 7'b0101100;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 7'b0101101;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 7'b0101110;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 7'b0101111;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 7'b0110000;
        state_var_NS = for_C_2;
      end
      for_C_2 : begin
        fsm_output = 7'b0110001;
        state_var_NS = for_C_3;
      end
      for_C_3 : begin
        fsm_output = 7'b0110010;
        state_var_NS = for_C_4;
      end
      for_C_4 : begin
        fsm_output = 7'b0110011;
        state_var_NS = for_C_5;
      end
      for_C_5 : begin
        fsm_output = 7'b0110100;
        state_var_NS = for_C_6;
      end
      for_C_6 : begin
        fsm_output = 7'b0110101;
        state_var_NS = for_C_7;
      end
      for_C_7 : begin
        fsm_output = 7'b0110110;
        state_var_NS = for_C_8;
      end
      for_C_8 : begin
        fsm_output = 7'b0110111;
        state_var_NS = for_C_9;
      end
      for_C_9 : begin
        fsm_output = 7'b0111000;
        state_var_NS = for_C_10;
      end
      for_C_10 : begin
        fsm_output = 7'b0111001;
        state_var_NS = for_C_11;
      end
      for_C_11 : begin
        fsm_output = 7'b0111010;
        state_var_NS = for_C_12;
      end
      for_C_12 : begin
        fsm_output = 7'b0111011;
        state_var_NS = for_C_13;
      end
      for_C_13 : begin
        fsm_output = 7'b0111100;
        state_var_NS = for_C_14;
      end
      for_C_14 : begin
        fsm_output = 7'b0111101;
        state_var_NS = for_C_15;
      end
      for_C_15 : begin
        fsm_output = 7'b0111110;
        state_var_NS = for_C_16;
      end
      for_C_16 : begin
        fsm_output = 7'b0111111;
        state_var_NS = for_C_17;
      end
      for_C_17 : begin
        fsm_output = 7'b1000000;
        state_var_NS = for_C_18;
      end
      for_C_18 : begin
        fsm_output = 7'b1000001;
        state_var_NS = for_C_19;
      end
      for_C_19 : begin
        fsm_output = 7'b1000010;
        state_var_NS = for_C_20;
      end
      for_C_20 : begin
        fsm_output = 7'b1000011;
        state_var_NS = for_C_21;
      end
      for_C_21 : begin
        fsm_output = 7'b1000100;
        state_var_NS = for_C_22;
      end
      for_C_22 : begin
        fsm_output = 7'b1000101;
        state_var_NS = for_C_23;
      end
      for_C_23 : begin
        fsm_output = 7'b1000110;
        state_var_NS = for_C_24;
      end
      for_C_24 : begin
        fsm_output = 7'b1000111;
        state_var_NS = for_C_25;
      end
      for_C_25 : begin
        fsm_output = 7'b1001000;
        state_var_NS = for_C_26;
      end
      for_C_26 : begin
        fsm_output = 7'b1001001;
        state_var_NS = for_C_27;
      end
      for_C_27 : begin
        fsm_output = 7'b1001010;
        state_var_NS = for_C_28;
      end
      for_C_28 : begin
        fsm_output = 7'b1001011;
        state_var_NS = for_C_29;
      end
      for_C_29 : begin
        fsm_output = 7'b1001100;
        state_var_NS = for_C_30;
      end
      for_C_30 : begin
        fsm_output = 7'b1001101;
        state_var_NS = for_C_31;
      end
      for_C_31 : begin
        fsm_output = 7'b1001110;
        state_var_NS = for_C_32;
      end
      for_C_32 : begin
        fsm_output = 7'b1001111;
        state_var_NS = for_C_33;
      end
      for_C_33 : begin
        fsm_output = 7'b1010000;
        state_var_NS = for_C_34;
      end
      for_C_34 : begin
        fsm_output = 7'b1010001;
        state_var_NS = for_C_35;
      end
      for_C_35 : begin
        fsm_output = 7'b1010010;
        state_var_NS = for_C_36;
      end
      for_C_36 : begin
        fsm_output = 7'b1010011;
        state_var_NS = for_C_37;
      end
      for_C_37 : begin
        fsm_output = 7'b1010100;
        state_var_NS = for_C_38;
      end
      for_C_38 : begin
        fsm_output = 7'b1010101;
        state_var_NS = for_C_39;
      end
      for_C_39 : begin
        fsm_output = 7'b1010110;
        state_var_NS = for_C_40;
      end
      for_C_40 : begin
        fsm_output = 7'b1010111;
        state_var_NS = for_C_41;
      end
      for_C_41 : begin
        fsm_output = 7'b1011000;
        if ( for_C_41_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 7'b0000000;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_staller
// ------------------------------------------------------------------


module ParamsDeserializer_run_staller (
  run_wen, inputChannel_rsci_wen_comp, qbuffer_params_rsci_wen_comp, render_params_rsci_wen_comp,
      accum_params_rsci_wen_comp, quad_serial_out_rsci_wen_comp
);
  output run_wen;
  input inputChannel_rsci_wen_comp;
  input qbuffer_params_rsci_wen_comp;
  input render_params_rsci_wen_comp;
  input accum_params_rsci_wen_comp;
  input quad_serial_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = inputChannel_rsci_wen_comp & qbuffer_params_rsci_wen_comp & render_params_rsci_wen_comp
      & accum_params_rsci_wen_comp & quad_serial_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_dp (
  clk, arst_n, quad_serial_out_rsci_oswt, quad_serial_out_rsci_wen_comp, quad_serial_out_rsci_biwt,
      quad_serial_out_rsci_bdwt, quad_serial_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_serial_out_rsci_oswt;
  output quad_serial_out_rsci_wen_comp;
  input quad_serial_out_rsci_biwt;
  input quad_serial_out_rsci_bdwt;
  output quad_serial_out_rsci_bcwt;
  reg quad_serial_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_serial_out_rsci_wen_comp = (~ quad_serial_out_rsci_oswt) | quad_serial_out_rsci_biwt
      | quad_serial_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_serial_out_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_serial_out_rsci_bcwt <= ~((~(quad_serial_out_rsci_bcwt | quad_serial_out_rsci_biwt))
          | quad_serial_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_ctrl (
  run_wen, quad_serial_out_rsci_oswt, quad_serial_out_rsci_irdy, quad_serial_out_rsci_biwt,
      quad_serial_out_rsci_bdwt, quad_serial_out_rsci_bcwt, quad_serial_out_rsci_ivld_run_sct
);
  input run_wen;
  input quad_serial_out_rsci_oswt;
  input quad_serial_out_rsci_irdy;
  output quad_serial_out_rsci_biwt;
  output quad_serial_out_rsci_bdwt;
  input quad_serial_out_rsci_bcwt;
  output quad_serial_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quad_serial_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_serial_out_rsci_bdwt = quad_serial_out_rsci_oswt & run_wen;
  assign quad_serial_out_rsci_biwt = quad_serial_out_rsci_ogwt & quad_serial_out_rsci_irdy;
  assign quad_serial_out_rsci_ogwt = quad_serial_out_rsci_oswt & (~ quad_serial_out_rsci_bcwt);
  assign quad_serial_out_rsci_ivld_run_sct = quad_serial_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_accum_params_rsci_accum_params_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_accum_params_rsci_accum_params_wait_dp (
  clk, arst_n, accum_params_rsci_oswt, accum_params_rsci_wen_comp, accum_params_rsci_biwt,
      accum_params_rsci_bdwt, accum_params_rsci_bcwt
);
  input clk;
  input arst_n;
  input accum_params_rsci_oswt;
  output accum_params_rsci_wen_comp;
  input accum_params_rsci_biwt;
  input accum_params_rsci_bdwt;
  output accum_params_rsci_bcwt;
  reg accum_params_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accum_params_rsci_wen_comp = (~ accum_params_rsci_oswt) | accum_params_rsci_biwt
      | accum_params_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accum_params_rsci_bcwt <= 1'b0;
    end
    else begin
      accum_params_rsci_bcwt <= ~((~(accum_params_rsci_bcwt | accum_params_rsci_biwt))
          | accum_params_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_accum_params_rsci_accum_params_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_accum_params_rsci_accum_params_wait_ctrl (
  run_wen, accum_params_rsci_oswt, accum_params_rsci_irdy, accum_params_rsci_biwt,
      accum_params_rsci_bdwt, accum_params_rsci_bcwt, accum_params_rsci_ivld_run_sct
);
  input run_wen;
  input accum_params_rsci_oswt;
  input accum_params_rsci_irdy;
  output accum_params_rsci_biwt;
  output accum_params_rsci_bdwt;
  input accum_params_rsci_bcwt;
  output accum_params_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire accum_params_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accum_params_rsci_bdwt = accum_params_rsci_oswt & run_wen;
  assign accum_params_rsci_biwt = accum_params_rsci_ogwt & accum_params_rsci_irdy;
  assign accum_params_rsci_ogwt = accum_params_rsci_oswt & (~ accum_params_rsci_bcwt);
  assign accum_params_rsci_ivld_run_sct = accum_params_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_render_params_rsci_render_params_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_render_params_rsci_render_params_wait_dp (
  clk, arst_n, render_params_rsci_oswt, render_params_rsci_wen_comp, render_params_rsci_biwt,
      render_params_rsci_bdwt, render_params_rsci_bcwt
);
  input clk;
  input arst_n;
  input render_params_rsci_oswt;
  output render_params_rsci_wen_comp;
  input render_params_rsci_biwt;
  input render_params_rsci_bdwt;
  output render_params_rsci_bcwt;
  reg render_params_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign render_params_rsci_wen_comp = (~ render_params_rsci_oswt) | render_params_rsci_biwt
      | render_params_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      render_params_rsci_bcwt <= 1'b0;
    end
    else begin
      render_params_rsci_bcwt <= ~((~(render_params_rsci_bcwt | render_params_rsci_biwt))
          | render_params_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_render_params_rsci_render_params_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_render_params_rsci_render_params_wait_ctrl (
  run_wen, render_params_rsci_oswt, render_params_rsci_irdy, render_params_rsci_biwt,
      render_params_rsci_bdwt, render_params_rsci_bcwt, render_params_rsci_ivld_run_sct
);
  input run_wen;
  input render_params_rsci_oswt;
  input render_params_rsci_irdy;
  output render_params_rsci_biwt;
  output render_params_rsci_bdwt;
  input render_params_rsci_bcwt;
  output render_params_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire render_params_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign render_params_rsci_bdwt = render_params_rsci_oswt & run_wen;
  assign render_params_rsci_biwt = render_params_rsci_ogwt & render_params_rsci_irdy;
  assign render_params_rsci_ogwt = render_params_rsci_oswt & (~ render_params_rsci_bcwt);
  assign render_params_rsci_ivld_run_sct = render_params_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_dp (
  clk, arst_n, qbuffer_params_rsci_oswt, qbuffer_params_rsci_wen_comp, qbuffer_params_rsci_biwt,
      qbuffer_params_rsci_bdwt, qbuffer_params_rsci_bcwt
);
  input clk;
  input arst_n;
  input qbuffer_params_rsci_oswt;
  output qbuffer_params_rsci_wen_comp;
  input qbuffer_params_rsci_biwt;
  input qbuffer_params_rsci_bdwt;
  output qbuffer_params_rsci_bcwt;
  reg qbuffer_params_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign qbuffer_params_rsci_wen_comp = (~ qbuffer_params_rsci_oswt) | qbuffer_params_rsci_biwt
      | qbuffer_params_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      qbuffer_params_rsci_bcwt <= 1'b0;
    end
    else begin
      qbuffer_params_rsci_bcwt <= ~((~(qbuffer_params_rsci_bcwt | qbuffer_params_rsci_biwt))
          | qbuffer_params_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_ctrl (
  run_wen, qbuffer_params_rsci_oswt, qbuffer_params_rsci_irdy, qbuffer_params_rsci_biwt,
      qbuffer_params_rsci_bdwt, qbuffer_params_rsci_bcwt, qbuffer_params_rsci_ivld_run_sct
);
  input run_wen;
  input qbuffer_params_rsci_oswt;
  input qbuffer_params_rsci_irdy;
  output qbuffer_params_rsci_biwt;
  output qbuffer_params_rsci_bdwt;
  input qbuffer_params_rsci_bcwt;
  output qbuffer_params_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire qbuffer_params_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign qbuffer_params_rsci_bdwt = qbuffer_params_rsci_oswt & run_wen;
  assign qbuffer_params_rsci_biwt = qbuffer_params_rsci_ogwt & qbuffer_params_rsci_irdy;
  assign qbuffer_params_rsci_ogwt = qbuffer_params_rsci_oswt & (~ qbuffer_params_rsci_bcwt);
  assign qbuffer_params_rsci_ivld_run_sct = qbuffer_params_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp (
  clk, arst_n, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt,
      inputChannel_rsci_biwt, inputChannel_rsci_bdwt, inputChannel_rsci_bcwt, inputChannel_rsci_idat
);
  input clk;
  input arst_n;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [11:0] inputChannel_rsci_idat_mxwt;
  input inputChannel_rsci_biwt;
  input inputChannel_rsci_bdwt;
  output inputChannel_rsci_bcwt;
  reg inputChannel_rsci_bcwt;
  input [11:0] inputChannel_rsci_idat;


  // Interconnect Declarations
  reg [11:0] inputChannel_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_wen_comp = (~ inputChannel_rsci_oswt) | inputChannel_rsci_biwt
      | inputChannel_rsci_bcwt;
  assign inputChannel_rsci_idat_mxwt = MUX_v_12_2_2(inputChannel_rsci_idat, inputChannel_rsci_idat_bfwt,
      inputChannel_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_bcwt <= 1'b0;
    end
    else begin
      inputChannel_rsci_bcwt <= ~((~(inputChannel_rsci_bcwt | inputChannel_rsci_biwt))
          | inputChannel_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_rsci_idat_bfwt <= 12'b000000000000;
    end
    else if ( ~ inputChannel_rsci_bcwt ) begin
      inputChannel_rsci_idat_bfwt <= inputChannel_rsci_idat_mxwt;
    end
  end

  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl (
  run_wen, inputChannel_rsci_oswt, inputChannel_rsci_biwt, inputChannel_rsci_bdwt,
      inputChannel_rsci_bcwt, inputChannel_rsci_irdy_run_sct, inputChannel_rsci_ivld
);
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_biwt;
  output inputChannel_rsci_bdwt;
  input inputChannel_rsci_bcwt;
  output inputChannel_rsci_irdy_run_sct;
  input inputChannel_rsci_ivld;


  // Interconnect Declarations
  wire inputChannel_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign inputChannel_rsci_bdwt = inputChannel_rsci_oswt & run_wen;
  assign inputChannel_rsci_biwt = inputChannel_rsci_ogwt & inputChannel_rsci_ivld;
  assign inputChannel_rsci_ogwt = inputChannel_rsci_oswt & (~ inputChannel_rsci_bcwt);
  assign inputChannel_rsci_irdy_run_sct = inputChannel_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_staller
// ------------------------------------------------------------------


module QuadBuffer_64_run_staller (
  run_wen, quads_in_rsci_wen_comp, paramsIn_rsci_wen_comp, quads_out_rsci_wen_comp
);
  output run_wen;
  input quads_in_rsci_wen_comp;
  input paramsIn_rsci_wen_comp;
  input quads_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = quads_in_rsci_wen_comp & paramsIn_rsci_wen_comp & quads_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_out_rsci_quads_out_wait_dp
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_out_rsci_quads_out_wait_dp (
  clk, arst_n, quads_out_rsci_oswt, quads_out_rsci_wen_comp, quads_out_rsci_biwt,
      quads_out_rsci_bdwt, quads_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input quads_out_rsci_oswt;
  output quads_out_rsci_wen_comp;
  input quads_out_rsci_biwt;
  input quads_out_rsci_bdwt;
  output quads_out_rsci_bcwt;
  reg quads_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quads_out_rsci_wen_comp = (~ quads_out_rsci_oswt) | quads_out_rsci_biwt
      | quads_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_out_rsci_bcwt <= 1'b0;
    end
    else begin
      quads_out_rsci_bcwt <= ~((~(quads_out_rsci_bcwt | quads_out_rsci_biwt)) | quads_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_out_rsci_quads_out_wait_ctrl
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_out_rsci_quads_out_wait_ctrl (
  run_wen, quads_out_rsci_oswt, quads_out_rsci_irdy, quads_out_rsci_biwt, quads_out_rsci_bdwt,
      quads_out_rsci_bcwt, quads_out_rsci_ivld_run_sct
);
  input run_wen;
  input quads_out_rsci_oswt;
  input quads_out_rsci_irdy;
  output quads_out_rsci_biwt;
  output quads_out_rsci_bdwt;
  input quads_out_rsci_bcwt;
  output quads_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quads_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_out_rsci_bdwt = quads_out_rsci_oswt & run_wen;
  assign quads_out_rsci_biwt = quads_out_rsci_ogwt & quads_out_rsci_irdy;
  assign quads_out_rsci_ogwt = quads_out_rsci_oswt & (~ quads_out_rsci_bcwt);
  assign quads_out_rsci_ivld_run_sct = quads_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [45:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [56:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  wire [56:0] paramsIn_rsci_idat_mxwt_pconst;
  reg [32:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [12:0] reg_paramsIn_rsci_idat_bfwt_ftd_12;
  reg reg_paramsIn_rsci_idat_bfwt_1_cse;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_pconst = MUX_v_57_2_2(paramsIn_rsci_idat, ({reg_paramsIn_rsci_idat_bfwt_ftd
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_ftd_12}),
      paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {(paramsIn_rsci_idat_mxwt_pconst[56:24]) , (paramsIn_rsci_idat_mxwt_pconst[12:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
      reg_paramsIn_rsci_idat_bfwt_1_cse <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
      reg_paramsIn_rsci_idat_bfwt_1_cse <= 1'b0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 33'b000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_pconst[56:24];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= 13'b0000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_12 <= paramsIn_rsci_idat_mxwt_pconst[12:0];
    end
  end

  function automatic [56:0] MUX_v_57_2_2;
    input [56:0] input_0;
    input [56:0] input_1;
    input [0:0] sel;
    reg [56:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_57_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_in_rsci_quads_in_wait_dp
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_in_rsci_quads_in_wait_dp (
  clk, arst_n, quads_in_rsci_oswt, quads_in_rsci_wen_comp, quads_in_rsci_idat_mxwt,
      quads_in_rsci_biwt, quads_in_rsci_bdwt, quads_in_rsci_bcwt, quads_in_rsci_idat
);
  input clk;
  input arst_n;
  input quads_in_rsci_oswt;
  output quads_in_rsci_wen_comp;
  output [376:0] quads_in_rsci_idat_mxwt;
  input quads_in_rsci_biwt;
  input quads_in_rsci_bdwt;
  output quads_in_rsci_bcwt;
  reg quads_in_rsci_bcwt;
  input [376:0] quads_in_rsci_idat;


  // Interconnect Declarations
  reg [376:0] quads_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_in_rsci_wen_comp = (~ quads_in_rsci_oswt) | quads_in_rsci_biwt | quads_in_rsci_bcwt;
  assign quads_in_rsci_idat_mxwt = MUX_v_377_2_2(quads_in_rsci_idat, quads_in_rsci_idat_bfwt,
      quads_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_in_rsci_bcwt <= 1'b0;
    end
    else begin
      quads_in_rsci_bcwt <= ~((~(quads_in_rsci_bcwt | quads_in_rsci_biwt)) | quads_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_in_rsci_idat_bfwt <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ quads_in_rsci_bcwt ) begin
      quads_in_rsci_idat_bfwt <= quads_in_rsci_idat_mxwt;
    end
  end

  function automatic [376:0] MUX_v_377_2_2;
    input [376:0] input_0;
    input [376:0] input_1;
    input [0:0] sel;
    reg [376:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_377_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_in_rsci_quads_in_wait_ctrl
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_in_rsci_quads_in_wait_ctrl (
  run_wen, quads_in_rsci_oswt, quads_in_rsci_biwt, quads_in_rsci_bdwt, quads_in_rsci_bcwt,
      quads_in_rsci_irdy_run_sct, quads_in_rsci_ivld
);
  input run_wen;
  input quads_in_rsci_oswt;
  output quads_in_rsci_biwt;
  output quads_in_rsci_bdwt;
  input quads_in_rsci_bcwt;
  output quads_in_rsci_irdy_run_sct;
  input quads_in_rsci_ivld;


  // Interconnect Declarations
  wire quads_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_in_rsci_bdwt = quads_in_rsci_oswt & run_wen;
  assign quads_in_rsci_biwt = quads_in_rsci_ogwt & quads_in_rsci_ivld;
  assign quads_in_rsci_ogwt = quads_in_rsci_oswt & (~ quads_in_rsci_bcwt);
  assign quads_in_rsci_irdy_run_sct = quads_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module RenderLooper_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for RenderLooper_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : RenderLooper_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_staller
// ------------------------------------------------------------------


module RenderLooper_run_staller (
  run_wen, render_params_rsci_wen_comp, render_params_out_rsci_wen_comp, loopIndicesOut_rsci_wen_comp
);
  output run_wen;
  input render_params_rsci_wen_comp;
  input render_params_out_rsci_wen_comp;
  input loopIndicesOut_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = render_params_rsci_wen_comp & render_params_out_rsci_wen_comp
      & loopIndicesOut_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp
// ------------------------------------------------------------------


module RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp (
  clk, arst_n, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input loopIndicesOut_rsci_biwt;
  input loopIndicesOut_rsci_bdwt;
  output loopIndicesOut_rsci_bcwt;
  reg loopIndicesOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_wen_comp = (~ loopIndicesOut_rsci_oswt) | loopIndicesOut_rsci_biwt
      | loopIndicesOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_bcwt <= 1'b0;
    end
    else begin
      loopIndicesOut_rsci_bcwt <= ~((~(loopIndicesOut_rsci_bcwt | loopIndicesOut_rsci_biwt))
          | loopIndicesOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl
// ------------------------------------------------------------------


module RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl (
  run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_irdy, loopIndicesOut_rsci_biwt,
      loopIndicesOut_rsci_bdwt, loopIndicesOut_rsci_bcwt, loopIndicesOut_rsci_ivld_run_sct
);
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  input loopIndicesOut_rsci_irdy;
  output loopIndicesOut_rsci_biwt;
  output loopIndicesOut_rsci_bdwt;
  input loopIndicesOut_rsci_bcwt;
  output loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesOut_rsci_bdwt = loopIndicesOut_rsci_oswt & run_wen;
  assign loopIndicesOut_rsci_biwt = loopIndicesOut_rsci_ogwt & loopIndicesOut_rsci_irdy;
  assign loopIndicesOut_rsci_ogwt = loopIndicesOut_rsci_oswt & (~ loopIndicesOut_rsci_bcwt);
  assign loopIndicesOut_rsci_ivld_run_sct = loopIndicesOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_out_rsci_render_params_out_wait_dp
// ------------------------------------------------------------------


module RenderLooper_run_render_params_out_rsci_render_params_out_wait_dp (
  clk, arst_n, render_params_out_rsci_oswt, render_params_out_rsci_wen_comp, render_params_out_rsci_biwt,
      render_params_out_rsci_bdwt, render_params_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input render_params_out_rsci_oswt;
  output render_params_out_rsci_wen_comp;
  input render_params_out_rsci_biwt;
  input render_params_out_rsci_bdwt;
  output render_params_out_rsci_bcwt;
  reg render_params_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign render_params_out_rsci_wen_comp = (~ render_params_out_rsci_oswt) | render_params_out_rsci_biwt
      | render_params_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      render_params_out_rsci_bcwt <= 1'b0;
    end
    else begin
      render_params_out_rsci_bcwt <= ~((~(render_params_out_rsci_bcwt | render_params_out_rsci_biwt))
          | render_params_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_out_rsci_render_params_out_wait_ctrl
// ------------------------------------------------------------------


module RenderLooper_run_render_params_out_rsci_render_params_out_wait_ctrl (
  run_wen, render_params_out_rsci_oswt, render_params_out_rsci_irdy, render_params_out_rsci_biwt,
      render_params_out_rsci_bdwt, render_params_out_rsci_bcwt, render_params_out_rsci_ivld_run_sct
);
  input run_wen;
  input render_params_out_rsci_oswt;
  input render_params_out_rsci_irdy;
  output render_params_out_rsci_biwt;
  output render_params_out_rsci_bdwt;
  input render_params_out_rsci_bcwt;
  output render_params_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire render_params_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign render_params_out_rsci_bdwt = render_params_out_rsci_oswt & run_wen;
  assign render_params_out_rsci_biwt = render_params_out_rsci_ogwt & render_params_out_rsci_irdy;
  assign render_params_out_rsci_ogwt = render_params_out_rsci_oswt & (~ render_params_out_rsci_bcwt);
  assign render_params_out_rsci_ivld_run_sct = render_params_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_rsci_render_params_wait_dp
// ------------------------------------------------------------------


module RenderLooper_run_render_params_rsci_render_params_wait_dp (
  clk, arst_n, render_params_rsci_oswt, render_params_rsci_wen_comp, render_params_rsci_idat_mxwt,
      render_params_rsci_biwt, render_params_rsci_bdwt, render_params_rsci_bcwt,
      render_params_rsci_idat
);
  input clk;
  input arst_n;
  input render_params_rsci_oswt;
  output render_params_rsci_wen_comp;
  output [419:0] render_params_rsci_idat_mxwt;
  input render_params_rsci_biwt;
  input render_params_rsci_bdwt;
  output render_params_rsci_bcwt;
  reg render_params_rsci_bcwt;
  input [419:0] render_params_rsci_idat;


  // Interconnect Declarations
  reg [419:0] render_params_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign render_params_rsci_wen_comp = (~ render_params_rsci_oswt) | render_params_rsci_biwt
      | render_params_rsci_bcwt;
  assign render_params_rsci_idat_mxwt = MUX_v_420_2_2(render_params_rsci_idat, render_params_rsci_idat_bfwt,
      render_params_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      render_params_rsci_bcwt <= 1'b0;
    end
    else begin
      render_params_rsci_bcwt <= ~((~(render_params_rsci_bcwt | render_params_rsci_biwt))
          | render_params_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      render_params_rsci_idat_bfwt <= 420'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ render_params_rsci_bcwt ) begin
      render_params_rsci_idat_bfwt <= render_params_rsci_idat_mxwt;
    end
  end

  function automatic [419:0] MUX_v_420_2_2;
    input [419:0] input_0;
    input [419:0] input_1;
    input [0:0] sel;
    reg [419:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_420_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_rsci_render_params_wait_ctrl
// ------------------------------------------------------------------


module RenderLooper_run_render_params_rsci_render_params_wait_ctrl (
  run_wen, render_params_rsci_oswt, render_params_rsci_biwt, render_params_rsci_bdwt,
      render_params_rsci_bcwt, render_params_rsci_irdy_run_sct, render_params_rsci_ivld
);
  input run_wen;
  input render_params_rsci_oswt;
  output render_params_rsci_biwt;
  output render_params_rsci_bdwt;
  input render_params_rsci_bcwt;
  output render_params_rsci_irdy_run_sct;
  input render_params_rsci_ivld;


  // Interconnect Declarations
  wire render_params_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign render_params_rsci_bdwt = render_params_rsci_oswt & run_wen;
  assign render_params_rsci_biwt = render_params_rsci_ogwt & render_params_rsci_ivld;
  assign render_params_rsci_ogwt = render_params_rsci_oswt & (~ render_params_rsci_bcwt);
  assign render_params_rsci_irdy_run_sct = render_params_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module RayGeneration_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for RayGeneration_run_run_fsm_1
  parameter
    run_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : RayGeneration_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_staller
// ------------------------------------------------------------------


module RayGeneration_run_staller (
  run_wen, loopIndicesIn_rsci_wen_comp, paramsIn_rsci_wen_comp, paramsOut_rsci_wen_comp,
      rayOut_rsci_wen_comp
);
  output run_wen;
  input loopIndicesIn_rsci_wen_comp;
  input paramsIn_rsci_wen_comp;
  input paramsOut_rsci_wen_comp;
  input rayOut_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = loopIndicesIn_rsci_wen_comp & paramsIn_rsci_wen_comp & paramsOut_rsci_wen_comp
      & rayOut_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_wait_dp
// ------------------------------------------------------------------


module RayGeneration_run_wait_dp (
  clk, arst_n, psq_vecMul1_run_mul_cmp_z, psq_vecMul1_run_mul_cmp_1_z, psq_vecMul1_run_mul_cmp_2_z,
      psq_vecMul1_run_mul_cmp_3_z, psq_vecMul1_run_mul_cmp_4_z, psq_vecMul1_run_mul_cmp_5_z,
      run_wen, psq_vecMul1_run_mul_cmp_z_oreg, psq_vecMul1_run_mul_cmp_1_z_oreg,
      psq_vecMul1_run_mul_cmp_2_z_oreg, psq_vecMul1_run_mul_cmp_3_z_oreg, psq_vecMul1_run_mul_cmp_4_z_oreg,
      psq_vecMul1_run_mul_cmp_5_z_oreg
);
  input clk;
  input arst_n;
  input [56:0] psq_vecMul1_run_mul_cmp_z;
  input [56:0] psq_vecMul1_run_mul_cmp_1_z;
  input [56:0] psq_vecMul1_run_mul_cmp_2_z;
  input [56:0] psq_vecMul1_run_mul_cmp_3_z;
  input [56:0] psq_vecMul1_run_mul_cmp_4_z;
  input [56:0] psq_vecMul1_run_mul_cmp_5_z;
  input run_wen;
  output [24:0] psq_vecMul1_run_mul_cmp_z_oreg;
  output [24:0] psq_vecMul1_run_mul_cmp_1_z_oreg;
  output [24:0] psq_vecMul1_run_mul_cmp_2_z_oreg;
  output [24:0] psq_vecMul1_run_mul_cmp_3_z_oreg;
  output [24:0] psq_vecMul1_run_mul_cmp_4_z_oreg;
  output [24:0] psq_vecMul1_run_mul_cmp_5_z_oreg;


  // Interconnect Declarations
  reg [24:0] psq_vecMul1_run_mul_cmp_z_oreg_pconst_56_32;
  reg [24:0] psq_vecMul1_run_mul_cmp_1_z_oreg_pconst_56_32;
  reg [24:0] psq_vecMul1_run_mul_cmp_2_z_oreg_pconst_56_32;
  reg [24:0] psq_vecMul1_run_mul_cmp_3_z_oreg_pconst_56_32;
  reg [24:0] psq_vecMul1_run_mul_cmp_4_z_oreg_pconst_56_32;
  reg [24:0] psq_vecMul1_run_mul_cmp_5_z_oreg_pconst_56_32;


  // Interconnect Declarations for Component Instantiations 
  assign psq_vecMul1_run_mul_cmp_z_oreg = psq_vecMul1_run_mul_cmp_z_oreg_pconst_56_32;
  assign psq_vecMul1_run_mul_cmp_1_z_oreg = psq_vecMul1_run_mul_cmp_1_z_oreg_pconst_56_32;
  assign psq_vecMul1_run_mul_cmp_2_z_oreg = psq_vecMul1_run_mul_cmp_2_z_oreg_pconst_56_32;
  assign psq_vecMul1_run_mul_cmp_3_z_oreg = psq_vecMul1_run_mul_cmp_3_z_oreg_pconst_56_32;
  assign psq_vecMul1_run_mul_cmp_4_z_oreg = psq_vecMul1_run_mul_cmp_4_z_oreg_pconst_56_32;
  assign psq_vecMul1_run_mul_cmp_5_z_oreg = psq_vecMul1_run_mul_cmp_5_z_oreg_pconst_56_32;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      psq_vecMul1_run_mul_cmp_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_1_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_2_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_3_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_4_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_5_z_oreg_pconst_56_32 <= 25'b0000000000000000000000000;
    end
    else if ( run_wen ) begin
      psq_vecMul1_run_mul_cmp_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_z[56:32];
      psq_vecMul1_run_mul_cmp_1_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_1_z[56:32];
      psq_vecMul1_run_mul_cmp_2_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_2_z[56:32];
      psq_vecMul1_run_mul_cmp_3_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_3_z[56:32];
      psq_vecMul1_run_mul_cmp_4_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_4_z[56:32];
      psq_vecMul1_run_mul_cmp_5_z_oreg_pconst_56_32 <= psq_vecMul1_run_mul_cmp_5_z[56:32];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_rayOut_rsci_rayOut_wait_dp
// ------------------------------------------------------------------


module RayGeneration_run_rayOut_rsci_rayOut_wait_dp (
  clk, arst_n, rayOut_rsci_oswt, rayOut_rsci_wen_comp, rayOut_rsci_biwt, rayOut_rsci_bdwt,
      rayOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input rayOut_rsci_oswt;
  output rayOut_rsci_wen_comp;
  input rayOut_rsci_biwt;
  input rayOut_rsci_bdwt;
  output rayOut_rsci_bcwt;
  reg rayOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rayOut_rsci_wen_comp = (~ rayOut_rsci_oswt) | rayOut_rsci_biwt | rayOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayOut_rsci_bcwt <= 1'b0;
    end
    else begin
      rayOut_rsci_bcwt <= ~((~(rayOut_rsci_bcwt | rayOut_rsci_biwt)) | rayOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_rayOut_rsci_rayOut_wait_ctrl
// ------------------------------------------------------------------


module RayGeneration_run_rayOut_rsci_rayOut_wait_ctrl (
  run_wen, rayOut_rsci_oswt, rayOut_rsci_irdy, rayOut_rsci_biwt, rayOut_rsci_bdwt,
      rayOut_rsci_bcwt, rayOut_rsci_ivld_run_sct
);
  input run_wen;
  input rayOut_rsci_oswt;
  input rayOut_rsci_irdy;
  output rayOut_rsci_biwt;
  output rayOut_rsci_bdwt;
  input rayOut_rsci_bcwt;
  output rayOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire rayOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rayOut_rsci_bdwt = rayOut_rsci_oswt & run_wen;
  assign rayOut_rsci_biwt = rayOut_rsci_ogwt & rayOut_rsci_irdy;
  assign rayOut_rsci_ogwt = rayOut_rsci_oswt & (~ rayOut_rsci_bcwt);
  assign rayOut_rsci_ivld_run_sct = rayOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsOut_rsci_paramsOut_wait_dp
// ------------------------------------------------------------------


module RayGeneration_run_paramsOut_rsci_paramsOut_wait_dp (
  clk, arst_n, paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_biwt,
      paramsOut_rsci_bdwt, paramsOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input paramsOut_rsci_biwt;
  input paramsOut_rsci_bdwt;
  output paramsOut_rsci_bcwt;
  reg paramsOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_wen_comp = (~ paramsOut_rsci_oswt) | paramsOut_rsci_biwt
      | paramsOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsOut_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsOut_rsci_bcwt <= ~((~(paramsOut_rsci_bcwt | paramsOut_rsci_biwt)) | paramsOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsOut_rsci_paramsOut_wait_ctrl
// ------------------------------------------------------------------


module RayGeneration_run_paramsOut_rsci_paramsOut_wait_ctrl (
  run_wen, paramsOut_rsci_oswt, paramsOut_rsci_irdy, paramsOut_rsci_biwt, paramsOut_rsci_bdwt,
      paramsOut_rsci_bcwt, paramsOut_rsci_ivld_run_sct
);
  input run_wen;
  input paramsOut_rsci_oswt;
  input paramsOut_rsci_irdy;
  output paramsOut_rsci_biwt;
  output paramsOut_rsci_bdwt;
  input paramsOut_rsci_bcwt;
  output paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire paramsOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_bdwt = paramsOut_rsci_oswt & run_wen;
  assign paramsOut_rsci_biwt = paramsOut_rsci_ogwt & paramsOut_rsci_irdy;
  assign paramsOut_rsci_ogwt = paramsOut_rsci_oswt & (~ paramsOut_rsci_bcwt);
  assign paramsOut_rsci_ivld_run_sct = paramsOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module RayGeneration_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [373:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [419:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  wire [419:0] paramsIn_rsci_idat_mxwt_pconst;
  reg [281:0] reg_paramsIn_rsci_idat_bfwt_ftd;
  reg [80:0] reg_paramsIn_rsci_idat_bfwt_ftd_45;
  reg [10:0] reg_paramsIn_rsci_idat_bfwt_ftd_48;
  reg reg_paramsIn_rsci_idat_bfwt_1_cse;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt_pconst = MUX_v_420_2_2(paramsIn_rsci_idat, ({reg_paramsIn_rsci_idat_bfwt_ftd
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_ftd_45
      , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_1_cse , reg_paramsIn_rsci_idat_bfwt_ftd_48}),
      paramsIn_rsci_bcwt);
  assign paramsIn_rsci_idat_mxwt = {(paramsIn_rsci_idat_mxwt_pconst[419:138]) , (paramsIn_rsci_idat_mxwt_pconst[93:13])
      , (paramsIn_rsci_idat_mxwt_pconst[10:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
      reg_paramsIn_rsci_idat_bfwt_1_cse <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
      reg_paramsIn_rsci_idat_bfwt_1_cse <= 1'b0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= 282'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd <= paramsIn_rsci_idat_mxwt_pconst[419:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_45 <= paramsIn_rsci_idat_mxwt_pconst[93:13];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_48 <= 11'b00000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      reg_paramsIn_rsci_idat_bfwt_ftd_48 <= paramsIn_rsci_idat_mxwt_pconst[10:0];
    end
  end

  function automatic [419:0] MUX_v_420_2_2;
    input [419:0] input_0;
    input [419:0] input_1;
    input [0:0] sel;
    reg [419:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_420_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module RayGeneration_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp
// ------------------------------------------------------------------


module RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp (
  clk, arst_n, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt,
      loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt, loopIndicesIn_rsci_bcwt,
      loopIndicesIn_rsci_idat
);
  input clk;
  input arst_n;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [22:0] loopIndicesIn_rsci_idat_mxwt;
  input loopIndicesIn_rsci_biwt;
  input loopIndicesIn_rsci_bdwt;
  output loopIndicesIn_rsci_bcwt;
  reg loopIndicesIn_rsci_bcwt;
  input [22:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations
  reg [22:0] loopIndicesIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_wen_comp = (~ loopIndicesIn_rsci_oswt) | loopIndicesIn_rsci_biwt
      | loopIndicesIn_rsci_bcwt;
  assign loopIndicesIn_rsci_idat_mxwt = MUX_v_23_2_2(loopIndicesIn_rsci_idat, loopIndicesIn_rsci_idat_bfwt,
      loopIndicesIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_rsci_bcwt <= 1'b0;
    end
    else begin
      loopIndicesIn_rsci_bcwt <= ~((~(loopIndicesIn_rsci_bcwt | loopIndicesIn_rsci_biwt))
          | loopIndicesIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesIn_rsci_idat_bfwt <= 23'b00000000000000000000000;
    end
    else if ( ~ loopIndicesIn_rsci_bcwt ) begin
      loopIndicesIn_rsci_idat_bfwt <= loopIndicesIn_rsci_idat_mxwt;
    end
  end

  function automatic [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl
// ------------------------------------------------------------------


module RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl (
  run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_biwt, loopIndicesIn_rsci_bdwt,
      loopIndicesIn_rsci_bcwt, loopIndicesIn_rsci_irdy_run_sct, loopIndicesIn_rsci_ivld
);
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_biwt;
  output loopIndicesIn_rsci_bdwt;
  input loopIndicesIn_rsci_bcwt;
  output loopIndicesIn_rsci_irdy_run_sct;
  input loopIndicesIn_rsci_ivld;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign loopIndicesIn_rsci_bdwt = loopIndicesIn_rsci_oswt & run_wen;
  assign loopIndicesIn_rsci_biwt = loopIndicesIn_rsci_ogwt & loopIndicesIn_rsci_ivld;
  assign loopIndicesIn_rsci_ogwt = loopIndicesIn_rsci_oswt & (~ loopIndicesIn_rsci_bcwt);
  assign loopIndicesIn_rsci_irdy_run_sct = loopIndicesIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module LoopDistrib_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, for_C_1_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input for_C_1_tr0;


  // FSM State Type Declaration for LoopDistrib_run_run_fsm_1
  parameter
    run_rlp_C_0 = 4'd0,
    main_C_0 = 4'd1,
    main_C_1 = 4'd2,
    main_C_2 = 4'd3,
    main_C_3 = 4'd4,
    main_C_4 = 4'd5,
    for_C_0 = 4'd6,
    for_C_1 = 4'd7,
    main_C_5 = 4'd8,
    main_C_6 = 4'd9;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : LoopDistrib_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 10'b0010000000;
        if ( for_C_1_tr0 ) begin
          state_var_NS = main_C_5;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_5 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 10'b0000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_staller
// ------------------------------------------------------------------


module LoopDistrib_run_staller (
  run_wen, ray_in_rsci_wen_comp, params_in_rsci_wen_comp, quads_rsci_wen_comp, attenuation_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_wen_comp, attenuation_chan_out_rsci_wen_comp,
      accumalated_color_out_rsci_wen_comp, ray_out_loopone_rsci_wen_comp, ray_out_looptwo_rsci_wen_comp,
      ray_out_worldhit_rsci_wen_comp, quad_out_loopone_rsci_wen_comp, quad_out_looptwo_rsci_wen_comp,
      quad_max_outone_rsci_wen_comp, quad_max_outtwo_rsci_wen_comp, params_out_rsci_wen_comp
);
  output run_wen;
  input ray_in_rsci_wen_comp;
  input params_in_rsci_wen_comp;
  input quads_rsci_wen_comp;
  input attenuation_chan_in_rsci_wen_comp;
  input accumalated_color_chan_in_rsci_wen_comp;
  input attenuation_chan_out_rsci_wen_comp;
  input accumalated_color_out_rsci_wen_comp;
  input ray_out_loopone_rsci_wen_comp;
  input ray_out_looptwo_rsci_wen_comp;
  input ray_out_worldhit_rsci_wen_comp;
  input quad_out_loopone_rsci_wen_comp;
  input quad_out_looptwo_rsci_wen_comp;
  input quad_max_outone_rsci_wen_comp;
  input quad_max_outtwo_rsci_wen_comp;
  input params_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = ray_in_rsci_wen_comp & params_in_rsci_wen_comp & quads_rsci_wen_comp
      & attenuation_chan_in_rsci_wen_comp & accumalated_color_chan_in_rsci_wen_comp
      & attenuation_chan_out_rsci_wen_comp & accumalated_color_out_rsci_wen_comp
      & ray_out_loopone_rsci_wen_comp & ray_out_looptwo_rsci_wen_comp & ray_out_worldhit_rsci_wen_comp
      & quad_out_loopone_rsci_wen_comp & quad_out_looptwo_rsci_wen_comp & quad_max_outone_rsci_wen_comp
      & quad_max_outtwo_rsci_wen_comp & params_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_out_rsci_params_out_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_params_out_rsci_params_out_wait_dp (
  clk, arst_n, params_out_rsci_oswt, params_out_rsci_wen_comp, params_out_rsci_biwt,
      params_out_rsci_bdwt, params_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input params_out_rsci_oswt;
  output params_out_rsci_wen_comp;
  input params_out_rsci_biwt;
  input params_out_rsci_bdwt;
  output params_out_rsci_bcwt;
  reg params_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign params_out_rsci_wen_comp = (~ params_out_rsci_oswt) | params_out_rsci_biwt
      | params_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_out_rsci_bcwt <= 1'b0;
    end
    else begin
      params_out_rsci_bcwt <= ~((~(params_out_rsci_bcwt | params_out_rsci_biwt))
          | params_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_out_rsci_params_out_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_params_out_rsci_params_out_wait_ctrl (
  run_wen, params_out_rsci_oswt, params_out_rsci_irdy, params_out_rsci_biwt, params_out_rsci_bdwt,
      params_out_rsci_bcwt, params_out_rsci_ivld_run_sct
);
  input run_wen;
  input params_out_rsci_oswt;
  input params_out_rsci_irdy;
  output params_out_rsci_biwt;
  output params_out_rsci_bdwt;
  input params_out_rsci_bcwt;
  output params_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire params_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_out_rsci_bdwt = params_out_rsci_oswt & run_wen;
  assign params_out_rsci_biwt = params_out_rsci_ogwt & params_out_rsci_irdy;
  assign params_out_rsci_ogwt = params_out_rsci_oswt & (~ params_out_rsci_bcwt);
  assign params_out_rsci_ivld_run_sct = params_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_dp (
  clk, arst_n, quad_max_outtwo_rsci_oswt, quad_max_outtwo_rsci_wen_comp, quad_max_outtwo_rsci_biwt,
      quad_max_outtwo_rsci_bdwt, quad_max_outtwo_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_max_outtwo_rsci_oswt;
  output quad_max_outtwo_rsci_wen_comp;
  input quad_max_outtwo_rsci_biwt;
  input quad_max_outtwo_rsci_bdwt;
  output quad_max_outtwo_rsci_bcwt;
  reg quad_max_outtwo_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_max_outtwo_rsci_wen_comp = (~ quad_max_outtwo_rsci_oswt) | quad_max_outtwo_rsci_biwt
      | quad_max_outtwo_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_outtwo_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_max_outtwo_rsci_bcwt <= ~((~(quad_max_outtwo_rsci_bcwt | quad_max_outtwo_rsci_biwt))
          | quad_max_outtwo_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_ctrl (
  run_wen, quad_max_outtwo_rsci_oswt, quad_max_outtwo_rsci_irdy, quad_max_outtwo_rsci_biwt,
      quad_max_outtwo_rsci_bdwt, quad_max_outtwo_rsci_bcwt, quad_max_outtwo_rsci_ivld_run_sct
);
  input run_wen;
  input quad_max_outtwo_rsci_oswt;
  input quad_max_outtwo_rsci_irdy;
  output quad_max_outtwo_rsci_biwt;
  output quad_max_outtwo_rsci_bdwt;
  input quad_max_outtwo_rsci_bcwt;
  output quad_max_outtwo_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quad_max_outtwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_max_outtwo_rsci_bdwt = quad_max_outtwo_rsci_oswt & run_wen;
  assign quad_max_outtwo_rsci_biwt = quad_max_outtwo_rsci_ogwt & quad_max_outtwo_rsci_irdy;
  assign quad_max_outtwo_rsci_ogwt = quad_max_outtwo_rsci_oswt & (~ quad_max_outtwo_rsci_bcwt);
  assign quad_max_outtwo_rsci_ivld_run_sct = quad_max_outtwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_dp (
  clk, arst_n, quad_max_outone_rsci_oswt, quad_max_outone_rsci_wen_comp, quad_max_outone_rsci_biwt,
      quad_max_outone_rsci_bdwt, quad_max_outone_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_max_outone_rsci_oswt;
  output quad_max_outone_rsci_wen_comp;
  input quad_max_outone_rsci_biwt;
  input quad_max_outone_rsci_bdwt;
  output quad_max_outone_rsci_bcwt;
  reg quad_max_outone_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_max_outone_rsci_wen_comp = (~ quad_max_outone_rsci_oswt) | quad_max_outone_rsci_biwt
      | quad_max_outone_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_outone_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_max_outone_rsci_bcwt <= ~((~(quad_max_outone_rsci_bcwt | quad_max_outone_rsci_biwt))
          | quad_max_outone_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_ctrl (
  run_wen, quad_max_outone_rsci_oswt, quad_max_outone_rsci_irdy, quad_max_outone_rsci_biwt,
      quad_max_outone_rsci_bdwt, quad_max_outone_rsci_bcwt, quad_max_outone_rsci_ivld_run_sct
);
  input run_wen;
  input quad_max_outone_rsci_oswt;
  input quad_max_outone_rsci_irdy;
  output quad_max_outone_rsci_biwt;
  output quad_max_outone_rsci_bdwt;
  input quad_max_outone_rsci_bcwt;
  output quad_max_outone_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quad_max_outone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_max_outone_rsci_bdwt = quad_max_outone_rsci_oswt & run_wen;
  assign quad_max_outone_rsci_biwt = quad_max_outone_rsci_ogwt & quad_max_outone_rsci_irdy;
  assign quad_max_outone_rsci_ogwt = quad_max_outone_rsci_oswt & (~ quad_max_outone_rsci_bcwt);
  assign quad_max_outone_rsci_ivld_run_sct = quad_max_outone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_dp (
  clk, arst_n, quad_out_looptwo_rsci_oswt, quad_out_looptwo_rsci_wen_comp, quad_out_looptwo_rsci_biwt,
      quad_out_looptwo_rsci_bdwt, quad_out_looptwo_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_out_looptwo_rsci_oswt;
  output quad_out_looptwo_rsci_wen_comp;
  input quad_out_looptwo_rsci_biwt;
  input quad_out_looptwo_rsci_bdwt;
  output quad_out_looptwo_rsci_bcwt;
  reg quad_out_looptwo_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_out_looptwo_rsci_wen_comp = (~ quad_out_looptwo_rsci_oswt) | quad_out_looptwo_rsci_biwt
      | quad_out_looptwo_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_out_looptwo_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_out_looptwo_rsci_bcwt <= ~((~(quad_out_looptwo_rsci_bcwt | quad_out_looptwo_rsci_biwt))
          | quad_out_looptwo_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_ctrl (
  run_wen, quad_out_looptwo_rsci_oswt, quad_out_looptwo_rsci_irdy, quad_out_looptwo_rsci_biwt,
      quad_out_looptwo_rsci_bdwt, quad_out_looptwo_rsci_bcwt, quad_out_looptwo_rsci_ivld_run_sct
);
  input run_wen;
  input quad_out_looptwo_rsci_oswt;
  input quad_out_looptwo_rsci_irdy;
  output quad_out_looptwo_rsci_biwt;
  output quad_out_looptwo_rsci_bdwt;
  input quad_out_looptwo_rsci_bcwt;
  output quad_out_looptwo_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quad_out_looptwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_out_looptwo_rsci_bdwt = quad_out_looptwo_rsci_oswt & run_wen;
  assign quad_out_looptwo_rsci_biwt = quad_out_looptwo_rsci_ogwt & quad_out_looptwo_rsci_irdy;
  assign quad_out_looptwo_rsci_ogwt = quad_out_looptwo_rsci_oswt & (~ quad_out_looptwo_rsci_bcwt);
  assign quad_out_looptwo_rsci_ivld_run_sct = quad_out_looptwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_dp (
  clk, arst_n, quad_out_loopone_rsci_oswt, quad_out_loopone_rsci_wen_comp, quad_out_loopone_rsci_biwt,
      quad_out_loopone_rsci_bdwt, quad_out_loopone_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_out_loopone_rsci_oswt;
  output quad_out_loopone_rsci_wen_comp;
  input quad_out_loopone_rsci_biwt;
  input quad_out_loopone_rsci_bdwt;
  output quad_out_loopone_rsci_bcwt;
  reg quad_out_loopone_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_out_loopone_rsci_wen_comp = (~ quad_out_loopone_rsci_oswt) | quad_out_loopone_rsci_biwt
      | quad_out_loopone_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_out_loopone_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_out_loopone_rsci_bcwt <= ~((~(quad_out_loopone_rsci_bcwt | quad_out_loopone_rsci_biwt))
          | quad_out_loopone_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_ctrl (
  run_wen, quad_out_loopone_rsci_oswt, quad_out_loopone_rsci_irdy, quad_out_loopone_rsci_biwt,
      quad_out_loopone_rsci_bdwt, quad_out_loopone_rsci_bcwt, quad_out_loopone_rsci_ivld_run_sct
);
  input run_wen;
  input quad_out_loopone_rsci_oswt;
  input quad_out_loopone_rsci_irdy;
  output quad_out_loopone_rsci_biwt;
  output quad_out_loopone_rsci_bdwt;
  input quad_out_loopone_rsci_bcwt;
  output quad_out_loopone_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire quad_out_loopone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_out_loopone_rsci_bdwt = quad_out_loopone_rsci_oswt & run_wen;
  assign quad_out_loopone_rsci_biwt = quad_out_loopone_rsci_ogwt & quad_out_loopone_rsci_irdy;
  assign quad_out_loopone_rsci_ogwt = quad_out_loopone_rsci_oswt & (~ quad_out_loopone_rsci_bcwt);
  assign quad_out_loopone_rsci_ivld_run_sct = quad_out_loopone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_dp (
  clk, arst_n, ray_out_worldhit_rsci_oswt, ray_out_worldhit_rsci_wen_comp, ray_out_worldhit_rsci_biwt,
      ray_out_worldhit_rsci_bdwt, ray_out_worldhit_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_worldhit_rsci_oswt;
  output ray_out_worldhit_rsci_wen_comp;
  input ray_out_worldhit_rsci_biwt;
  input ray_out_worldhit_rsci_bdwt;
  output ray_out_worldhit_rsci_bcwt;
  reg ray_out_worldhit_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_worldhit_rsci_wen_comp = (~ ray_out_worldhit_rsci_oswt) | ray_out_worldhit_rsci_biwt
      | ray_out_worldhit_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_worldhit_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_worldhit_rsci_bcwt <= ~((~(ray_out_worldhit_rsci_bcwt | ray_out_worldhit_rsci_biwt))
          | ray_out_worldhit_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_ctrl (
  run_wen, ray_out_worldhit_rsci_oswt, ray_out_worldhit_rsci_irdy, ray_out_worldhit_rsci_biwt,
      ray_out_worldhit_rsci_bdwt, ray_out_worldhit_rsci_bcwt, ray_out_worldhit_rsci_ivld_run_sct
);
  input run_wen;
  input ray_out_worldhit_rsci_oswt;
  input ray_out_worldhit_rsci_irdy;
  output ray_out_worldhit_rsci_biwt;
  output ray_out_worldhit_rsci_bdwt;
  input ray_out_worldhit_rsci_bcwt;
  output ray_out_worldhit_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire ray_out_worldhit_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_worldhit_rsci_bdwt = ray_out_worldhit_rsci_oswt & run_wen;
  assign ray_out_worldhit_rsci_biwt = ray_out_worldhit_rsci_ogwt & ray_out_worldhit_rsci_irdy;
  assign ray_out_worldhit_rsci_ogwt = ray_out_worldhit_rsci_oswt & (~ ray_out_worldhit_rsci_bcwt);
  assign ray_out_worldhit_rsci_ivld_run_sct = ray_out_worldhit_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_dp (
  clk, arst_n, ray_out_looptwo_rsci_oswt, ray_out_looptwo_rsci_wen_comp, ray_out_looptwo_rsci_biwt,
      ray_out_looptwo_rsci_bdwt, ray_out_looptwo_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_looptwo_rsci_oswt;
  output ray_out_looptwo_rsci_wen_comp;
  input ray_out_looptwo_rsci_biwt;
  input ray_out_looptwo_rsci_bdwt;
  output ray_out_looptwo_rsci_bcwt;
  reg ray_out_looptwo_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_looptwo_rsci_wen_comp = (~ ray_out_looptwo_rsci_oswt) | ray_out_looptwo_rsci_biwt
      | ray_out_looptwo_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_looptwo_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_looptwo_rsci_bcwt <= ~((~(ray_out_looptwo_rsci_bcwt | ray_out_looptwo_rsci_biwt))
          | ray_out_looptwo_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_ctrl (
  run_wen, ray_out_looptwo_rsci_oswt, ray_out_looptwo_rsci_irdy, ray_out_looptwo_rsci_biwt,
      ray_out_looptwo_rsci_bdwt, ray_out_looptwo_rsci_bcwt, ray_out_looptwo_rsci_ivld_run_sct
);
  input run_wen;
  input ray_out_looptwo_rsci_oswt;
  input ray_out_looptwo_rsci_irdy;
  output ray_out_looptwo_rsci_biwt;
  output ray_out_looptwo_rsci_bdwt;
  input ray_out_looptwo_rsci_bcwt;
  output ray_out_looptwo_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire ray_out_looptwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_looptwo_rsci_bdwt = ray_out_looptwo_rsci_oswt & run_wen;
  assign ray_out_looptwo_rsci_biwt = ray_out_looptwo_rsci_ogwt & ray_out_looptwo_rsci_irdy;
  assign ray_out_looptwo_rsci_ogwt = ray_out_looptwo_rsci_oswt & (~ ray_out_looptwo_rsci_bcwt);
  assign ray_out_looptwo_rsci_ivld_run_sct = ray_out_looptwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_dp (
  clk, arst_n, ray_out_loopone_rsci_oswt, ray_out_loopone_rsci_wen_comp, ray_out_loopone_rsci_biwt,
      ray_out_loopone_rsci_bdwt, ray_out_loopone_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_loopone_rsci_oswt;
  output ray_out_loopone_rsci_wen_comp;
  input ray_out_loopone_rsci_biwt;
  input ray_out_loopone_rsci_bdwt;
  output ray_out_loopone_rsci_bcwt;
  reg ray_out_loopone_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_loopone_rsci_wen_comp = (~ ray_out_loopone_rsci_oswt) | ray_out_loopone_rsci_biwt
      | ray_out_loopone_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_loopone_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_loopone_rsci_bcwt <= ~((~(ray_out_loopone_rsci_bcwt | ray_out_loopone_rsci_biwt))
          | ray_out_loopone_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_ctrl (
  run_wen, ray_out_loopone_rsci_oswt, ray_out_loopone_rsci_irdy, ray_out_loopone_rsci_biwt,
      ray_out_loopone_rsci_bdwt, ray_out_loopone_rsci_bcwt, ray_out_loopone_rsci_ivld_run_sct
);
  input run_wen;
  input ray_out_loopone_rsci_oswt;
  input ray_out_loopone_rsci_irdy;
  output ray_out_loopone_rsci_biwt;
  output ray_out_loopone_rsci_bdwt;
  input ray_out_loopone_rsci_bcwt;
  output ray_out_loopone_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire ray_out_loopone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_loopone_rsci_bdwt = ray_out_loopone_rsci_oswt & run_wen;
  assign ray_out_loopone_rsci_biwt = ray_out_loopone_rsci_ogwt & ray_out_loopone_rsci_irdy;
  assign ray_out_loopone_rsci_ogwt = ray_out_loopone_rsci_oswt & (~ ray_out_loopone_rsci_bcwt);
  assign ray_out_loopone_rsci_ivld_run_sct = ray_out_loopone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_dp (
  clk, arst_n, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_biwt, accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input accumalated_color_out_rsci_biwt;
  input accumalated_color_out_rsci_bdwt;
  output accumalated_color_out_rsci_bcwt;
  reg accumalated_color_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_wen_comp = (~ accumalated_color_out_rsci_oswt)
      | accumalated_color_out_rsci_biwt | accumalated_color_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_out_rsci_bcwt <= ~((~(accumalated_color_out_rsci_bcwt | accumalated_color_out_rsci_biwt))
          | accumalated_color_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
    (
  run_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_irdy, accumalated_color_out_rsci_biwt,
      accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt, accumalated_color_out_rsci_ivld_run_sct
);
  input run_wen;
  input accumalated_color_out_rsci_oswt;
  input accumalated_color_out_rsci_irdy;
  output accumalated_color_out_rsci_biwt;
  output accumalated_color_out_rsci_bdwt;
  input accumalated_color_out_rsci_bcwt;
  output accumalated_color_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_bdwt = accumalated_color_out_rsci_oswt & run_wen;
  assign accumalated_color_out_rsci_biwt = accumalated_color_out_rsci_ogwt & accumalated_color_out_rsci_irdy;
  assign accumalated_color_out_rsci_ogwt = accumalated_color_out_rsci_oswt & (~ accumalated_color_out_rsci_bcwt);
  assign accumalated_color_out_rsci_ivld_run_sct = accumalated_color_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp (
  clk, arst_n, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_biwt, attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input attenuation_chan_out_rsci_biwt;
  input attenuation_chan_out_rsci_bdwt;
  output attenuation_chan_out_rsci_bcwt;
  reg attenuation_chan_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_wen_comp = (~ attenuation_chan_out_rsci_oswt)
      | attenuation_chan_out_rsci_biwt | attenuation_chan_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_out_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_out_rsci_bcwt <= ~((~(attenuation_chan_out_rsci_bcwt | attenuation_chan_out_rsci_biwt))
          | attenuation_chan_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl (
  run_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_irdy, attenuation_chan_out_rsci_biwt,
      attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt, attenuation_chan_out_rsci_ivld_run_sct
);
  input run_wen;
  input attenuation_chan_out_rsci_oswt;
  input attenuation_chan_out_rsci_irdy;
  output attenuation_chan_out_rsci_biwt;
  output attenuation_chan_out_rsci_bdwt;
  input attenuation_chan_out_rsci_bcwt;
  output attenuation_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_bdwt = attenuation_chan_out_rsci_oswt & run_wen;
  assign attenuation_chan_out_rsci_biwt = attenuation_chan_out_rsci_ogwt & attenuation_chan_out_rsci_irdy;
  assign attenuation_chan_out_rsci_ogwt = attenuation_chan_out_rsci_oswt & (~ attenuation_chan_out_rsci_bcwt);
  assign attenuation_chan_out_rsci_ivld_run_sct = attenuation_chan_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
    (
  clk, arst_n, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_idat_mxwt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  input accumalated_color_chan_in_rsci_biwt;
  input accumalated_color_chan_in_rsci_bdwt;
  output accumalated_color_chan_in_rsci_bcwt;
  reg accumalated_color_chan_in_rsci_bcwt;
  input [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] accumalated_color_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_wen_comp = (~ accumalated_color_chan_in_rsci_oswt)
      | accumalated_color_chan_in_rsci_biwt | accumalated_color_chan_in_rsci_bcwt;
  assign accumalated_color_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(accumalated_color_chan_in_rsci_idat,
      accumalated_color_chan_in_rsci_idat_bfwt, accumalated_color_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_chan_in_rsci_bcwt <= ~((~(accumalated_color_chan_in_rsci_bcwt
          | accumalated_color_chan_in_rsci_biwt)) | accumalated_color_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ accumalated_color_chan_in_rsci_bcwt ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
    (
  run_wen, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_irdy_run_sct,
      accumalated_color_chan_in_rsci_ivld
);
  input run_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_biwt;
  output accumalated_color_chan_in_rsci_bdwt;
  input accumalated_color_chan_in_rsci_bcwt;
  output accumalated_color_chan_in_rsci_irdy_run_sct;
  input accumalated_color_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_bdwt = accumalated_color_chan_in_rsci_oswt
      & run_wen;
  assign accumalated_color_chan_in_rsci_biwt = accumalated_color_chan_in_rsci_ogwt
      & accumalated_color_chan_in_rsci_ivld;
  assign accumalated_color_chan_in_rsci_ogwt = accumalated_color_chan_in_rsci_oswt
      & (~ accumalated_color_chan_in_rsci_bcwt);
  assign accumalated_color_chan_in_rsci_irdy_run_sct = accumalated_color_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp (
  clk, arst_n, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;
  input attenuation_chan_in_rsci_biwt;
  input attenuation_chan_in_rsci_bdwt;
  output attenuation_chan_in_rsci_bcwt;
  reg attenuation_chan_in_rsci_bcwt;
  input [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] attenuation_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_wen_comp = (~ attenuation_chan_in_rsci_oswt) |
      attenuation_chan_in_rsci_biwt | attenuation_chan_in_rsci_bcwt;
  assign attenuation_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(attenuation_chan_in_rsci_idat,
      attenuation_chan_in_rsci_idat_bfwt, attenuation_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_in_rsci_bcwt <= ~((~(attenuation_chan_in_rsci_bcwt | attenuation_chan_in_rsci_biwt))
          | attenuation_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ attenuation_chan_in_rsci_bcwt ) begin
      attenuation_chan_in_rsci_idat_bfwt <= attenuation_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl (
  run_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_irdy_run_sct, attenuation_chan_in_rsci_ivld
);
  input run_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_biwt;
  output attenuation_chan_in_rsci_bdwt;
  input attenuation_chan_in_rsci_bcwt;
  output attenuation_chan_in_rsci_irdy_run_sct;
  input attenuation_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_bdwt = attenuation_chan_in_rsci_oswt & run_wen;
  assign attenuation_chan_in_rsci_biwt = attenuation_chan_in_rsci_ogwt & attenuation_chan_in_rsci_ivld;
  assign attenuation_chan_in_rsci_ogwt = attenuation_chan_in_rsci_oswt & (~ attenuation_chan_in_rsci_bcwt);
  assign attenuation_chan_in_rsci_irdy_run_sct = attenuation_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quads_rsci_quads_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_quads_rsci_quads_wait_dp (
  clk, arst_n, quads_rsci_oswt, quads_rsci_wen_comp, quads_rsci_idat_mxwt, quads_rsci_biwt,
      quads_rsci_bdwt, quads_rsci_bcwt, quads_rsci_idat
);
  input clk;
  input arst_n;
  input quads_rsci_oswt;
  output quads_rsci_wen_comp;
  output [376:0] quads_rsci_idat_mxwt;
  input quads_rsci_biwt;
  input quads_rsci_bdwt;
  output quads_rsci_bcwt;
  reg quads_rsci_bcwt;
  input [376:0] quads_rsci_idat;


  // Interconnect Declarations
  reg [376:0] quads_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_rsci_wen_comp = (~ quads_rsci_oswt) | quads_rsci_biwt | quads_rsci_bcwt;
  assign quads_rsci_idat_mxwt = MUX_v_377_2_2(quads_rsci_idat, quads_rsci_idat_bfwt,
      quads_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_rsci_bcwt <= 1'b0;
    end
    else begin
      quads_rsci_bcwt <= ~((~(quads_rsci_bcwt | quads_rsci_biwt)) | quads_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_rsci_idat_bfwt <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ quads_rsci_bcwt ) begin
      quads_rsci_idat_bfwt <= quads_rsci_idat_mxwt;
    end
  end

  function automatic [376:0] MUX_v_377_2_2;
    input [376:0] input_0;
    input [376:0] input_1;
    input [0:0] sel;
    reg [376:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_377_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quads_rsci_quads_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_quads_rsci_quads_wait_ctrl (
  run_wen, quads_rsci_oswt, quads_rsci_biwt, quads_rsci_bdwt, quads_rsci_bcwt, quads_rsci_irdy_run_sct,
      quads_rsci_ivld
);
  input run_wen;
  input quads_rsci_oswt;
  output quads_rsci_biwt;
  output quads_rsci_bdwt;
  input quads_rsci_bcwt;
  output quads_rsci_irdy_run_sct;
  input quads_rsci_ivld;


  // Interconnect Declarations
  wire quads_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_rsci_bdwt = quads_rsci_oswt & run_wen;
  assign quads_rsci_biwt = quads_rsci_ogwt & quads_rsci_ivld;
  assign quads_rsci_ogwt = quads_rsci_oswt & (~ quads_rsci_bcwt);
  assign quads_rsci_irdy_run_sct = quads_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_in_rsci_params_in_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_params_in_rsci_params_in_wait_dp (
  clk, arst_n, params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt,
      params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt, params_in_rsci_idat
);
  input clk;
  input arst_n;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [92:0] params_in_rsci_idat_mxwt;
  input params_in_rsci_biwt;
  input params_in_rsci_bdwt;
  output params_in_rsci_bcwt;
  reg params_in_rsci_bcwt;
  input [92:0] params_in_rsci_idat;


  // Interconnect Declarations
  reg [92:0] params_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_wen_comp = (~ params_in_rsci_oswt) | params_in_rsci_biwt
      | params_in_rsci_bcwt;
  assign params_in_rsci_idat_mxwt = MUX_v_93_2_2(params_in_rsci_idat, params_in_rsci_idat_bfwt,
      params_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_bcwt <= 1'b0;
    end
    else begin
      params_in_rsci_bcwt <= ~((~(params_in_rsci_bcwt | params_in_rsci_biwt)) | params_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_idat_bfwt <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ params_in_rsci_bcwt ) begin
      params_in_rsci_idat_bfwt <= params_in_rsci_idat_mxwt;
    end
  end

  function automatic [92:0] MUX_v_93_2_2;
    input [92:0] input_0;
    input [92:0] input_1;
    input [0:0] sel;
    reg [92:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_93_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_in_rsci_params_in_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_params_in_rsci_params_in_wait_ctrl (
  run_wen, params_in_rsci_oswt, params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt,
      params_in_rsci_irdy_run_sct, params_in_rsci_ivld
);
  input run_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_biwt;
  output params_in_rsci_bdwt;
  input params_in_rsci_bcwt;
  output params_in_rsci_irdy_run_sct;
  input params_in_rsci_ivld;


  // Interconnect Declarations
  wire params_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_bdwt = params_in_rsci_oswt & run_wen;
  assign params_in_rsci_biwt = params_in_rsci_ogwt & params_in_rsci_ivld;
  assign params_in_rsci_ogwt = params_in_rsci_oswt & (~ params_in_rsci_bcwt);
  assign params_in_rsci_irdy_run_sct = params_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_in_rsci_ray_in_wait_dp
// ------------------------------------------------------------------


module LoopDistrib_run_ray_in_rsci_ray_in_wait_dp (
  clk, arst_n, ray_in_rsci_oswt, ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt, ray_in_rsci_biwt,
      ray_in_rsci_bdwt, ray_in_rsci_bcwt, ray_in_rsci_idat
);
  input clk;
  input arst_n;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [165:0] ray_in_rsci_idat_mxwt;
  input ray_in_rsci_biwt;
  input ray_in_rsci_bdwt;
  output ray_in_rsci_bcwt;
  reg ray_in_rsci_bcwt;
  input [165:0] ray_in_rsci_idat;


  // Interconnect Declarations
  reg [165:0] ray_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_wen_comp = (~ ray_in_rsci_oswt) | ray_in_rsci_biwt | ray_in_rsci_bcwt;
  assign ray_in_rsci_idat_mxwt = MUX_v_166_2_2(ray_in_rsci_idat, ray_in_rsci_idat_bfwt,
      ray_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_in_rsci_bcwt <= ~((~(ray_in_rsci_bcwt | ray_in_rsci_biwt)) | ray_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_in_rsci_bcwt ) begin
      ray_in_rsci_idat_bfwt <= ray_in_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_in_rsci_ray_in_wait_ctrl
// ------------------------------------------------------------------


module LoopDistrib_run_ray_in_rsci_ray_in_wait_ctrl (
  run_wen, ray_in_rsci_oswt, ray_in_rsci_biwt, ray_in_rsci_bdwt, ray_in_rsci_bcwt,
      ray_in_rsci_irdy_run_sct, ray_in_rsci_ivld
);
  input run_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_biwt;
  output ray_in_rsci_bdwt;
  input ray_in_rsci_bcwt;
  output ray_in_rsci_irdy_run_sct;
  input ray_in_rsci_ivld;


  // Interconnect Declarations
  wire ray_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_bdwt = ray_in_rsci_oswt & run_wen;
  assign ray_in_rsci_biwt = ray_in_rsci_ogwt & ray_in_rsci_ivld;
  assign ray_in_rsci_ogwt = ray_in_rsci_oswt & (~ ray_in_rsci_bcwt);
  assign ray_in_rsci_irdy_run_sct = ray_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_hit_fsm
//  FSM Module
// ------------------------------------------------------------------


module IntersecLoop_hit_hit_fsm (
  clk, arst_n, hit_wen, fsm_output, for_C_3_tr0
);
  input clk;
  input arst_n;
  input hit_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input for_C_3_tr0;


  // FSM State Type Declaration for IntersecLoop_hit_hit_fsm_1
  parameter
    hit_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    for_C_0 = 3'd2,
    for_C_1 = 3'd3,
    for_C_2 = 3'd4,
    for_C_3 = 3'd5,
    main_C_1 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : IntersecLoop_hit_hit_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 7'b0000010;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 7'b0000100;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 7'b0001000;
        state_var_NS = for_C_2;
      end
      for_C_2 : begin
        fsm_output = 7'b0010000;
        state_var_NS = for_C_3;
      end
      for_C_3 : begin
        fsm_output = 7'b0100000;
        if ( for_C_3_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // hit_rlp_C_0
      default : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= hit_rlp_C_0;
    end
    else if ( hit_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_staller
// ------------------------------------------------------------------


module IntersecLoop_hit_staller (
  hit_wen, quads_rsci_wen_comp, ray_temp_in_rsci_wen_comp, quad_max_in_rsci_wen_comp,
      quad_hit_anything_out_rsci_wen_comp, rec_quad_out_rsci_wen_comp, closest_so_far_out_rsci_wen_comp
);
  output hit_wen;
  input quads_rsci_wen_comp;
  input ray_temp_in_rsci_wen_comp;
  input quad_max_in_rsci_wen_comp;
  input quad_hit_anything_out_rsci_wen_comp;
  input rec_quad_out_rsci_wen_comp;
  input closest_so_far_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign hit_wen = quads_rsci_wen_comp & ray_temp_in_rsci_wen_comp & quad_max_in_rsci_wen_comp
      & quad_hit_anything_out_rsci_wen_comp & rec_quad_out_rsci_wen_comp & closest_so_far_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_wait_dp (
  clk, arst_n, ensig_cgo_iro, mult_run_mul_cmp_en, mult_run_mul_cmp_z, quadInters_qnorm_rorig_run_mul_1_cmp_z,
      quadInters_qnorm_rorig_run_mul_1_cmp_1_z, quadInters_qnorm_rorig_run_mul_1_cmp_2_z,
      quadInters_qnorm_rorig_run_mul_1_cmp_3_z, quadInters_qnorm_rorig_run_mul_1_cmp_4_z,
      quadInters_qnorm_rorig_run_mul_1_cmp_5_z, quadInters_denom_dot_run_mul_2_cmp_z,
      quadInters_denom_dot_run_mul_2_cmp_1_z, quadInters_denom_dot_run_mul_1_cmp_z,
      hit_wen, ensig_cgo, mult_run_mul_cmp_z_oreg, quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg,
      quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg, quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg,
      quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg, quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg,
      quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg, quadInters_denom_dot_run_mul_2_cmp_z_oreg,
      quadInters_denom_dot_run_mul_2_cmp_1_z_oreg, quadInters_denom_dot_run_mul_1_cmp_z_oreg
);
  input clk;
  input arst_n;
  input ensig_cgo_iro;
  output mult_run_mul_cmp_en;
  input [74:0] mult_run_mul_cmp_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_z;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_z;
  input [57:0] quadInters_denom_dot_run_mul_2_cmp_z;
  input [57:0] quadInters_denom_dot_run_mul_2_cmp_1_z;
  input [59:0] quadInters_denom_dot_run_mul_1_cmp_z;
  input hit_wen;
  input ensig_cgo;
  output [44:0] mult_run_mul_cmp_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg;
  output [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg;
  reg [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg;
  output [57:0] quadInters_denom_dot_run_mul_2_cmp_z_oreg;
  reg [57:0] quadInters_denom_dot_run_mul_2_cmp_z_oreg;
  output [57:0] quadInters_denom_dot_run_mul_2_cmp_1_z_oreg;
  reg [57:0] quadInters_denom_dot_run_mul_2_cmp_1_z_oreg;
  output [59:0] quadInters_denom_dot_run_mul_1_cmp_z_oreg;
  reg [59:0] quadInters_denom_dot_run_mul_1_cmp_z_oreg;


  // Interconnect Declarations
  reg [44:0] mult_run_mul_cmp_z_oreg_pconst_74_30;


  // Interconnect Declarations for Component Instantiations 
  assign mult_run_mul_cmp_en = ~(hit_wen & (ensig_cgo | ensig_cgo_iro));
  assign mult_run_mul_cmp_z_oreg = mult_run_mul_cmp_z_oreg_pconst_74_30;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mult_run_mul_cmp_z_oreg_pconst_74_30 <= 45'b000000000000000000000000000000000000000000000;
    end
    else if ( ~ mult_run_mul_cmp_en ) begin
      mult_run_mul_cmp_z_oreg_pconst_74_30 <= mult_run_mul_cmp_z[74:30];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg <= 62'b00000000000000000000000000000000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_z_oreg <= 58'b0000000000000000000000000000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_1_z_oreg <= 58'b0000000000000000000000000000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_1_cmp_z_oreg <= 60'b000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( hit_wen ) begin
      quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_z;
      quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_1_z;
      quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_2_z;
      quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_3_z;
      quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_4_z;
      quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg <= quadInters_qnorm_rorig_run_mul_1_cmp_5_z;
      quadInters_denom_dot_run_mul_2_cmp_z_oreg <= quadInters_denom_dot_run_mul_2_cmp_z;
      quadInters_denom_dot_run_mul_2_cmp_1_z_oreg <= quadInters_denom_dot_run_mul_2_cmp_1_z;
      quadInters_denom_dot_run_mul_1_cmp_z_oreg <= quadInters_denom_dot_run_mul_1_cmp_z;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_dp (
  clk, arst_n, closest_so_far_out_rsci_oswt, closest_so_far_out_rsci_wen_comp, closest_so_far_out_rsci_biwt,
      closest_so_far_out_rsci_bdwt, closest_so_far_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input closest_so_far_out_rsci_oswt;
  output closest_so_far_out_rsci_wen_comp;
  input closest_so_far_out_rsci_biwt;
  input closest_so_far_out_rsci_bdwt;
  output closest_so_far_out_rsci_bcwt;
  reg closest_so_far_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_out_rsci_wen_comp = (~ closest_so_far_out_rsci_oswt) | closest_so_far_out_rsci_biwt
      | closest_so_far_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_out_rsci_bcwt <= 1'b0;
    end
    else begin
      closest_so_far_out_rsci_bcwt <= ~((~(closest_so_far_out_rsci_bcwt | closest_so_far_out_rsci_biwt))
          | closest_so_far_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_ctrl (
  hit_wen, closest_so_far_out_rsci_oswt, closest_so_far_out_rsci_irdy, closest_so_far_out_rsci_biwt,
      closest_so_far_out_rsci_bdwt, closest_so_far_out_rsci_bcwt, closest_so_far_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input closest_so_far_out_rsci_oswt;
  input closest_so_far_out_rsci_irdy;
  output closest_so_far_out_rsci_biwt;
  output closest_so_far_out_rsci_bdwt;
  input closest_so_far_out_rsci_bcwt;
  output closest_so_far_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire closest_so_far_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_out_rsci_bdwt = closest_so_far_out_rsci_oswt & hit_wen;
  assign closest_so_far_out_rsci_biwt = closest_so_far_out_rsci_ogwt & closest_so_far_out_rsci_irdy;
  assign closest_so_far_out_rsci_ogwt = closest_so_far_out_rsci_oswt & (~ closest_so_far_out_rsci_bcwt);
  assign closest_so_far_out_rsci_ivld_hit_sct = closest_so_far_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_dp (
  clk, arst_n, rec_quad_out_rsci_oswt, rec_quad_out_rsci_wen_comp, rec_quad_out_rsci_biwt,
      rec_quad_out_rsci_bdwt, rec_quad_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input rec_quad_out_rsci_oswt;
  output rec_quad_out_rsci_wen_comp;
  input rec_quad_out_rsci_biwt;
  input rec_quad_out_rsci_bdwt;
  output rec_quad_out_rsci_bcwt;
  reg rec_quad_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_out_rsci_wen_comp = (~ rec_quad_out_rsci_oswt) | rec_quad_out_rsci_biwt
      | rec_quad_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_out_rsci_bcwt <= 1'b0;
    end
    else begin
      rec_quad_out_rsci_bcwt <= ~((~(rec_quad_out_rsci_bcwt | rec_quad_out_rsci_biwt))
          | rec_quad_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_ctrl (
  hit_wen, rec_quad_out_rsci_oswt, rec_quad_out_rsci_irdy, rec_quad_out_rsci_biwt,
      rec_quad_out_rsci_bdwt, rec_quad_out_rsci_bcwt, rec_quad_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input rec_quad_out_rsci_oswt;
  input rec_quad_out_rsci_irdy;
  output rec_quad_out_rsci_biwt;
  output rec_quad_out_rsci_bdwt;
  input rec_quad_out_rsci_bcwt;
  output rec_quad_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire rec_quad_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_out_rsci_bdwt = rec_quad_out_rsci_oswt & hit_wen;
  assign rec_quad_out_rsci_biwt = rec_quad_out_rsci_ogwt & rec_quad_out_rsci_irdy;
  assign rec_quad_out_rsci_ogwt = rec_quad_out_rsci_oswt & (~ rec_quad_out_rsci_bcwt);
  assign rec_quad_out_rsci_ivld_hit_sct = rec_quad_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_dp
    (
  clk, arst_n, quad_hit_anything_out_rsci_oswt, quad_hit_anything_out_rsci_wen_comp,
      quad_hit_anything_out_rsci_biwt, quad_hit_anything_out_rsci_bdwt, quad_hit_anything_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input quad_hit_anything_out_rsci_oswt;
  output quad_hit_anything_out_rsci_wen_comp;
  input quad_hit_anything_out_rsci_biwt;
  input quad_hit_anything_out_rsci_bdwt;
  output quad_hit_anything_out_rsci_bcwt;
  reg quad_hit_anything_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_out_rsci_wen_comp = (~ quad_hit_anything_out_rsci_oswt)
      | quad_hit_anything_out_rsci_biwt | quad_hit_anything_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_out_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_hit_anything_out_rsci_bcwt <= ~((~(quad_hit_anything_out_rsci_bcwt | quad_hit_anything_out_rsci_biwt))
          | quad_hit_anything_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_ctrl
    (
  hit_wen, quad_hit_anything_out_rsci_oswt, quad_hit_anything_out_rsci_irdy, quad_hit_anything_out_rsci_biwt,
      quad_hit_anything_out_rsci_bdwt, quad_hit_anything_out_rsci_bcwt, quad_hit_anything_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input quad_hit_anything_out_rsci_oswt;
  input quad_hit_anything_out_rsci_irdy;
  output quad_hit_anything_out_rsci_biwt;
  output quad_hit_anything_out_rsci_bdwt;
  input quad_hit_anything_out_rsci_bcwt;
  output quad_hit_anything_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire quad_hit_anything_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_out_rsci_bdwt = quad_hit_anything_out_rsci_oswt & hit_wen;
  assign quad_hit_anything_out_rsci_biwt = quad_hit_anything_out_rsci_ogwt & quad_hit_anything_out_rsci_irdy;
  assign quad_hit_anything_out_rsci_ogwt = quad_hit_anything_out_rsci_oswt & (~ quad_hit_anything_out_rsci_bcwt);
  assign quad_hit_anything_out_rsci_ivld_hit_sct = quad_hit_anything_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_dp (
  clk, arst_n, quad_max_in_rsci_oswt, quad_max_in_rsci_wen_comp, quad_max_in_rsci_idat_mxwt,
      quad_max_in_rsci_biwt, quad_max_in_rsci_bdwt, quad_max_in_rsci_bcwt, quad_max_in_rsci_idat
);
  input clk;
  input arst_n;
  input quad_max_in_rsci_oswt;
  output quad_max_in_rsci_wen_comp;
  output [10:0] quad_max_in_rsci_idat_mxwt;
  input quad_max_in_rsci_biwt;
  input quad_max_in_rsci_bdwt;
  output quad_max_in_rsci_bcwt;
  reg quad_max_in_rsci_bcwt;
  input [10:0] quad_max_in_rsci_idat;


  // Interconnect Declarations
  reg [10:0] quad_max_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_max_in_rsci_wen_comp = (~ quad_max_in_rsci_oswt) | quad_max_in_rsci_biwt
      | quad_max_in_rsci_bcwt;
  assign quad_max_in_rsci_idat_mxwt = MUX_v_11_2_2(quad_max_in_rsci_idat, quad_max_in_rsci_idat_bfwt,
      quad_max_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_in_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_max_in_rsci_bcwt <= ~((~(quad_max_in_rsci_bcwt | quad_max_in_rsci_biwt))
          | quad_max_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_in_rsci_idat_bfwt <= 11'b00000000000;
    end
    else if ( ~ quad_max_in_rsci_bcwt ) begin
      quad_max_in_rsci_idat_bfwt <= quad_max_in_rsci_idat_mxwt;
    end
  end

  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_ctrl (
  hit_wen, quad_max_in_rsci_oswt, quad_max_in_rsci_biwt, quad_max_in_rsci_bdwt, quad_max_in_rsci_bcwt,
      quad_max_in_rsci_irdy_hit_sct, quad_max_in_rsci_ivld
);
  input hit_wen;
  input quad_max_in_rsci_oswt;
  output quad_max_in_rsci_biwt;
  output quad_max_in_rsci_bdwt;
  input quad_max_in_rsci_bcwt;
  output quad_max_in_rsci_irdy_hit_sct;
  input quad_max_in_rsci_ivld;


  // Interconnect Declarations
  wire quad_max_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_max_in_rsci_bdwt = quad_max_in_rsci_oswt & hit_wen;
  assign quad_max_in_rsci_biwt = quad_max_in_rsci_ogwt & quad_max_in_rsci_ivld;
  assign quad_max_in_rsci_ogwt = quad_max_in_rsci_oswt & (~ quad_max_in_rsci_bcwt);
  assign quad_max_in_rsci_irdy_hit_sct = quad_max_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_dp (
  clk, arst_n, ray_temp_in_rsci_oswt, ray_temp_in_rsci_wen_comp, ray_temp_in_rsci_idat_mxwt,
      ray_temp_in_rsci_biwt, ray_temp_in_rsci_bdwt, ray_temp_in_rsci_bcwt, ray_temp_in_rsci_idat
);
  input clk;
  input arst_n;
  input ray_temp_in_rsci_oswt;
  output ray_temp_in_rsci_wen_comp;
  output [165:0] ray_temp_in_rsci_idat_mxwt;
  input ray_temp_in_rsci_biwt;
  input ray_temp_in_rsci_bdwt;
  output ray_temp_in_rsci_bcwt;
  reg ray_temp_in_rsci_bcwt;
  input [165:0] ray_temp_in_rsci_idat;


  // Interconnect Declarations
  reg [165:0] ray_temp_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_temp_in_rsci_wen_comp = (~ ray_temp_in_rsci_oswt) | ray_temp_in_rsci_biwt
      | ray_temp_in_rsci_bcwt;
  assign ray_temp_in_rsci_idat_mxwt = MUX_v_166_2_2(ray_temp_in_rsci_idat, ray_temp_in_rsci_idat_bfwt,
      ray_temp_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_temp_in_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_temp_in_rsci_bcwt <= ~((~(ray_temp_in_rsci_bcwt | ray_temp_in_rsci_biwt))
          | ray_temp_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_temp_in_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_temp_in_rsci_bcwt ) begin
      ray_temp_in_rsci_idat_bfwt <= ray_temp_in_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_ctrl (
  hit_wen, ray_temp_in_rsci_oswt, ray_temp_in_rsci_biwt, ray_temp_in_rsci_bdwt, ray_temp_in_rsci_bcwt,
      ray_temp_in_rsci_irdy_hit_sct, ray_temp_in_rsci_ivld
);
  input hit_wen;
  input ray_temp_in_rsci_oswt;
  output ray_temp_in_rsci_biwt;
  output ray_temp_in_rsci_bdwt;
  input ray_temp_in_rsci_bcwt;
  output ray_temp_in_rsci_irdy_hit_sct;
  input ray_temp_in_rsci_ivld;


  // Interconnect Declarations
  wire ray_temp_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_temp_in_rsci_bdwt = ray_temp_in_rsci_oswt & hit_wen;
  assign ray_temp_in_rsci_biwt = ray_temp_in_rsci_ogwt & ray_temp_in_rsci_ivld;
  assign ray_temp_in_rsci_ogwt = ray_temp_in_rsci_oswt & (~ ray_temp_in_rsci_bcwt);
  assign ray_temp_in_rsci_irdy_hit_sct = ray_temp_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quads_rsci_quads_wait_dp
// ------------------------------------------------------------------


module IntersecLoop_hit_quads_rsci_quads_wait_dp (
  clk, arst_n, quads_rsci_oswt, quads_rsci_wen_comp, quads_rsci_idat_mxwt, quads_rsci_biwt,
      quads_rsci_bdwt, quads_rsci_bcwt, quads_rsci_idat
);
  input clk;
  input arst_n;
  input quads_rsci_oswt;
  output quads_rsci_wen_comp;
  output [376:0] quads_rsci_idat_mxwt;
  input quads_rsci_biwt;
  input quads_rsci_bdwt;
  output quads_rsci_bcwt;
  reg quads_rsci_bcwt;
  input [376:0] quads_rsci_idat;


  // Interconnect Declarations
  reg [376:0] quads_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_rsci_wen_comp = (~ quads_rsci_oswt) | quads_rsci_biwt | quads_rsci_bcwt;
  assign quads_rsci_idat_mxwt = MUX_v_377_2_2(quads_rsci_idat, quads_rsci_idat_bfwt,
      quads_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_rsci_bcwt <= 1'b0;
    end
    else begin
      quads_rsci_bcwt <= ~((~(quads_rsci_bcwt | quads_rsci_biwt)) | quads_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_rsci_idat_bfwt <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ quads_rsci_bcwt ) begin
      quads_rsci_idat_bfwt <= quads_rsci_idat_mxwt;
    end
  end

  function automatic [376:0] MUX_v_377_2_2;
    input [376:0] input_0;
    input [376:0] input_1;
    input [0:0] sel;
    reg [376:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_377_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quads_rsci_quads_wait_ctrl
// ------------------------------------------------------------------


module IntersecLoop_hit_quads_rsci_quads_wait_ctrl (
  hit_wen, quads_rsci_oswt, quads_rsci_biwt, quads_rsci_bdwt, quads_rsci_bcwt, quads_rsci_irdy_hit_sct,
      quads_rsci_ivld
);
  input hit_wen;
  input quads_rsci_oswt;
  output quads_rsci_biwt;
  output quads_rsci_bdwt;
  input quads_rsci_bcwt;
  output quads_rsci_irdy_hit_sct;
  input quads_rsci_ivld;


  // Interconnect Declarations
  wire quads_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quads_rsci_bdwt = quads_rsci_oswt & hit_wen;
  assign quads_rsci_biwt = quads_rsci_ogwt & quads_rsci_ivld;
  assign quads_rsci_ogwt = quads_rsci_oswt & (~ quads_rsci_bcwt);
  assign quads_rsci_irdy_hit_sct = quads_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_hit_fsm
//  FSM Module
// ------------------------------------------------------------------


module WorldHit_hit_hit_fsm (
  clk, arst_n, hit_wen, fsm_output
);
  input clk;
  input arst_n;
  input hit_wen;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;


  // FSM State Type Declaration for WorldHit_hit_hit_fsm_1
  parameter
    hit_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    main_C_1 = 3'd2,
    main_C_2 = 3'd3,
    main_C_3 = 3'd4,
    main_C_4 = 3'd5,
    main_C_5 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : WorldHit_hit_hit_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 7'b0000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 7'b0000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b0001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b0010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 7'b0100000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // hit_rlp_C_0
      default : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= hit_rlp_C_0;
    end
    else if ( hit_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_staller
// ------------------------------------------------------------------


module WorldHit_hit_staller (
  hit_wen, ray_in_rsci_wen_comp, params_in_rsci_wen_comp, attenuation_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_wen_comp, quad_hit_anything_outone_rsci_wen_comp,
      quad_hit_anything_outtwo_rsci_wen_comp, rec_quad_outone_rsci_wen_comp, rec_quad_outtwo_rsci_wen_comp,
      closest_so_far_outone_rsci_wen_comp, closest_so_far_outtwo_rsci_wen_comp, attenuation_chan_out_rsci_wen_comp,
      accumalated_color_out_rsci_wen_comp, hit_out_rsci_wen_comp, ray_out_rsci_wen_comp,
      isHit_rsci_wen_comp
);
  output hit_wen;
  input ray_in_rsci_wen_comp;
  input params_in_rsci_wen_comp;
  input attenuation_chan_in_rsci_wen_comp;
  input accumalated_color_chan_in_rsci_wen_comp;
  input quad_hit_anything_outone_rsci_wen_comp;
  input quad_hit_anything_outtwo_rsci_wen_comp;
  input rec_quad_outone_rsci_wen_comp;
  input rec_quad_outtwo_rsci_wen_comp;
  input closest_so_far_outone_rsci_wen_comp;
  input closest_so_far_outtwo_rsci_wen_comp;
  input attenuation_chan_out_rsci_wen_comp;
  input accumalated_color_out_rsci_wen_comp;
  input hit_out_rsci_wen_comp;
  input ray_out_rsci_wen_comp;
  input isHit_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign hit_wen = ray_in_rsci_wen_comp & params_in_rsci_wen_comp & attenuation_chan_in_rsci_wen_comp
      & accumalated_color_chan_in_rsci_wen_comp & quad_hit_anything_outone_rsci_wen_comp
      & quad_hit_anything_outtwo_rsci_wen_comp & rec_quad_outone_rsci_wen_comp &
      rec_quad_outtwo_rsci_wen_comp & closest_so_far_outone_rsci_wen_comp & closest_so_far_outtwo_rsci_wen_comp
      & attenuation_chan_out_rsci_wen_comp & accumalated_color_out_rsci_wen_comp
      & hit_out_rsci_wen_comp & ray_out_rsci_wen_comp & isHit_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_wait_dp (
  clk, arst_n, else_mul_cmp_z, hit_wen, else_mul_cmp_z_oreg
);
  input clk;
  input arst_n;
  input [48:0] else_mul_cmp_z;
  input hit_wen;
  output [26:0] else_mul_cmp_z_oreg;


  // Interconnect Declarations
  reg [26:0] else_mul_cmp_z_oreg_pconst_48_22;


  // Interconnect Declarations for Component Instantiations 
  assign else_mul_cmp_z_oreg = else_mul_cmp_z_oreg_pconst_48_22;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      else_mul_cmp_z_oreg_pconst_48_22 <= 27'b000000000000000000000000000;
    end
    else if ( hit_wen ) begin
      else_mul_cmp_z_oreg_pconst_48_22 <= else_mul_cmp_z[48:22];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_isHit_rsci_isHit_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_isHit_rsci_isHit_wait_dp (
  clk, arst_n, isHit_rsci_oswt, isHit_rsci_wen_comp, isHit_rsci_biwt, isHit_rsci_bdwt,
      isHit_rsci_bcwt
);
  input clk;
  input arst_n;
  input isHit_rsci_oswt;
  output isHit_rsci_wen_comp;
  input isHit_rsci_biwt;
  input isHit_rsci_bdwt;
  output isHit_rsci_bcwt;
  reg isHit_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign isHit_rsci_wen_comp = (~ isHit_rsci_oswt) | isHit_rsci_biwt | isHit_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      isHit_rsci_bcwt <= 1'b0;
    end
    else begin
      isHit_rsci_bcwt <= ~((~(isHit_rsci_bcwt | isHit_rsci_biwt)) | isHit_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_isHit_rsci_isHit_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_isHit_rsci_isHit_wait_ctrl (
  hit_wen, isHit_rsci_oswt, isHit_rsci_irdy, isHit_rsci_biwt, isHit_rsci_bdwt, isHit_rsci_bcwt,
      isHit_rsci_ivld_hit_sct
);
  input hit_wen;
  input isHit_rsci_oswt;
  input isHit_rsci_irdy;
  output isHit_rsci_biwt;
  output isHit_rsci_bdwt;
  input isHit_rsci_bcwt;
  output isHit_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire isHit_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign isHit_rsci_bdwt = isHit_rsci_oswt & hit_wen;
  assign isHit_rsci_biwt = isHit_rsci_ogwt & isHit_rsci_irdy;
  assign isHit_rsci_ogwt = isHit_rsci_oswt & (~ isHit_rsci_bcwt);
  assign isHit_rsci_ivld_hit_sct = isHit_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_out_rsci_ray_out_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_ray_out_rsci_ray_out_wait_dp (
  clk, arst_n, ray_out_rsci_oswt, ray_out_rsci_wen_comp, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input ray_out_rsci_biwt;
  input ray_out_rsci_bdwt;
  output ray_out_rsci_bcwt;
  reg ray_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_wen_comp = (~ ray_out_rsci_oswt) | ray_out_rsci_biwt | ray_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_rsci_bcwt <= ~((~(ray_out_rsci_bcwt | ray_out_rsci_biwt)) | ray_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_out_rsci_ray_out_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_ray_out_rsci_ray_out_wait_ctrl (
  hit_wen, ray_out_rsci_oswt, ray_out_rsci_irdy, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt, ray_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input ray_out_rsci_oswt;
  input ray_out_rsci_irdy;
  output ray_out_rsci_biwt;
  output ray_out_rsci_bdwt;
  input ray_out_rsci_bcwt;
  output ray_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire ray_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_bdwt = ray_out_rsci_oswt & hit_wen;
  assign ray_out_rsci_biwt = ray_out_rsci_ogwt & ray_out_rsci_irdy;
  assign ray_out_rsci_ogwt = ray_out_rsci_oswt & (~ ray_out_rsci_bcwt);
  assign ray_out_rsci_ivld_hit_sct = ray_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_hit_out_rsci_hit_out_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_hit_out_rsci_hit_out_wait_dp (
  clk, arst_n, hit_out_rsci_oswt, hit_out_rsci_wen_comp, hit_out_rsci_biwt, hit_out_rsci_bdwt,
      hit_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input hit_out_rsci_oswt;
  output hit_out_rsci_wen_comp;
  input hit_out_rsci_biwt;
  input hit_out_rsci_bdwt;
  output hit_out_rsci_bcwt;
  reg hit_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign hit_out_rsci_wen_comp = (~ hit_out_rsci_oswt) | hit_out_rsci_biwt | hit_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      hit_out_rsci_bcwt <= 1'b0;
    end
    else begin
      hit_out_rsci_bcwt <= ~((~(hit_out_rsci_bcwt | hit_out_rsci_biwt)) | hit_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_hit_out_rsci_hit_out_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_hit_out_rsci_hit_out_wait_ctrl (
  hit_wen, hit_out_rsci_oswt, hit_out_rsci_irdy, hit_out_rsci_biwt, hit_out_rsci_bdwt,
      hit_out_rsci_bcwt, hit_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input hit_out_rsci_oswt;
  input hit_out_rsci_irdy;
  output hit_out_rsci_biwt;
  output hit_out_rsci_bdwt;
  input hit_out_rsci_bcwt;
  output hit_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire hit_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign hit_out_rsci_bdwt = hit_out_rsci_oswt & hit_wen;
  assign hit_out_rsci_biwt = hit_out_rsci_ogwt & hit_out_rsci_irdy;
  assign hit_out_rsci_ogwt = hit_out_rsci_oswt & (~ hit_out_rsci_bcwt);
  assign hit_out_rsci_ivld_hit_sct = hit_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_dp (
  clk, arst_n, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_biwt, accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input accumalated_color_out_rsci_biwt;
  input accumalated_color_out_rsci_bdwt;
  output accumalated_color_out_rsci_bcwt;
  reg accumalated_color_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_wen_comp = (~ accumalated_color_out_rsci_oswt)
      | accumalated_color_out_rsci_biwt | accumalated_color_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_out_rsci_bcwt <= ~((~(accumalated_color_out_rsci_bcwt | accumalated_color_out_rsci_biwt))
          | accumalated_color_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl (
  hit_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_irdy, accumalated_color_out_rsci_biwt,
      accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt, accumalated_color_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input accumalated_color_out_rsci_oswt;
  input accumalated_color_out_rsci_irdy;
  output accumalated_color_out_rsci_biwt;
  output accumalated_color_out_rsci_bdwt;
  input accumalated_color_out_rsci_bcwt;
  output accumalated_color_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_bdwt = accumalated_color_out_rsci_oswt & hit_wen;
  assign accumalated_color_out_rsci_biwt = accumalated_color_out_rsci_ogwt & accumalated_color_out_rsci_irdy;
  assign accumalated_color_out_rsci_ogwt = accumalated_color_out_rsci_oswt & (~ accumalated_color_out_rsci_bcwt);
  assign accumalated_color_out_rsci_ivld_hit_sct = accumalated_color_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp (
  clk, arst_n, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_biwt, attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input attenuation_chan_out_rsci_biwt;
  input attenuation_chan_out_rsci_bdwt;
  output attenuation_chan_out_rsci_bcwt;
  reg attenuation_chan_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_wen_comp = (~ attenuation_chan_out_rsci_oswt)
      | attenuation_chan_out_rsci_biwt | attenuation_chan_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_out_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_out_rsci_bcwt <= ~((~(attenuation_chan_out_rsci_bcwt | attenuation_chan_out_rsci_biwt))
          | attenuation_chan_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl (
  hit_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_irdy, attenuation_chan_out_rsci_biwt,
      attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt, attenuation_chan_out_rsci_ivld_hit_sct
);
  input hit_wen;
  input attenuation_chan_out_rsci_oswt;
  input attenuation_chan_out_rsci_irdy;
  output attenuation_chan_out_rsci_biwt;
  output attenuation_chan_out_rsci_bdwt;
  input attenuation_chan_out_rsci_bcwt;
  output attenuation_chan_out_rsci_ivld_hit_sct;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_bdwt = attenuation_chan_out_rsci_oswt & hit_wen;
  assign attenuation_chan_out_rsci_biwt = attenuation_chan_out_rsci_ogwt & attenuation_chan_out_rsci_irdy;
  assign attenuation_chan_out_rsci_ogwt = attenuation_chan_out_rsci_oswt & (~ attenuation_chan_out_rsci_bcwt);
  assign attenuation_chan_out_rsci_ivld_hit_sct = attenuation_chan_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_dp (
  clk, arst_n, closest_so_far_outtwo_rsci_oswt, closest_so_far_outtwo_rsci_wen_comp,
      closest_so_far_outtwo_rsci_idat_mxwt, closest_so_far_outtwo_rsci_biwt, closest_so_far_outtwo_rsci_bdwt,
      closest_so_far_outtwo_rsci_bcwt, closest_so_far_outtwo_rsci_idat
);
  input clk;
  input arst_n;
  input closest_so_far_outtwo_rsci_oswt;
  output closest_so_far_outtwo_rsci_wen_comp;
  output [46:0] closest_so_far_outtwo_rsci_idat_mxwt;
  input closest_so_far_outtwo_rsci_biwt;
  input closest_so_far_outtwo_rsci_bdwt;
  output closest_so_far_outtwo_rsci_bcwt;
  reg closest_so_far_outtwo_rsci_bcwt;
  input [46:0] closest_so_far_outtwo_rsci_idat;


  // Interconnect Declarations
  reg [46:0] closest_so_far_outtwo_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_outtwo_rsci_wen_comp = (~ closest_so_far_outtwo_rsci_oswt)
      | closest_so_far_outtwo_rsci_biwt | closest_so_far_outtwo_rsci_bcwt;
  assign closest_so_far_outtwo_rsci_idat_mxwt = MUX_v_47_2_2(closest_so_far_outtwo_rsci_idat,
      closest_so_far_outtwo_rsci_idat_bfwt, closest_so_far_outtwo_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_outtwo_rsci_bcwt <= 1'b0;
    end
    else begin
      closest_so_far_outtwo_rsci_bcwt <= ~((~(closest_so_far_outtwo_rsci_bcwt | closest_so_far_outtwo_rsci_biwt))
          | closest_so_far_outtwo_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_outtwo_rsci_idat_bfwt <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( ~ closest_so_far_outtwo_rsci_bcwt ) begin
      closest_so_far_outtwo_rsci_idat_bfwt <= closest_so_far_outtwo_rsci_idat_mxwt;
    end
  end

  function automatic [46:0] MUX_v_47_2_2;
    input [46:0] input_0;
    input [46:0] input_1;
    input [0:0] sel;
    reg [46:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_47_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_ctrl (
  hit_wen, closest_so_far_outtwo_rsci_oswt, closest_so_far_outtwo_rsci_biwt, closest_so_far_outtwo_rsci_bdwt,
      closest_so_far_outtwo_rsci_bcwt, closest_so_far_outtwo_rsci_irdy_hit_sct, closest_so_far_outtwo_rsci_ivld
);
  input hit_wen;
  input closest_so_far_outtwo_rsci_oswt;
  output closest_so_far_outtwo_rsci_biwt;
  output closest_so_far_outtwo_rsci_bdwt;
  input closest_so_far_outtwo_rsci_bcwt;
  output closest_so_far_outtwo_rsci_irdy_hit_sct;
  input closest_so_far_outtwo_rsci_ivld;


  // Interconnect Declarations
  wire closest_so_far_outtwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_outtwo_rsci_bdwt = closest_so_far_outtwo_rsci_oswt & hit_wen;
  assign closest_so_far_outtwo_rsci_biwt = closest_so_far_outtwo_rsci_ogwt & closest_so_far_outtwo_rsci_ivld;
  assign closest_so_far_outtwo_rsci_ogwt = closest_so_far_outtwo_rsci_oswt & (~ closest_so_far_outtwo_rsci_bcwt);
  assign closest_so_far_outtwo_rsci_irdy_hit_sct = closest_so_far_outtwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_dp (
  clk, arst_n, closest_so_far_outone_rsci_oswt, closest_so_far_outone_rsci_wen_comp,
      closest_so_far_outone_rsci_idat_mxwt, closest_so_far_outone_rsci_biwt, closest_so_far_outone_rsci_bdwt,
      closest_so_far_outone_rsci_bcwt, closest_so_far_outone_rsci_idat
);
  input clk;
  input arst_n;
  input closest_so_far_outone_rsci_oswt;
  output closest_so_far_outone_rsci_wen_comp;
  output [46:0] closest_so_far_outone_rsci_idat_mxwt;
  input closest_so_far_outone_rsci_biwt;
  input closest_so_far_outone_rsci_bdwt;
  output closest_so_far_outone_rsci_bcwt;
  reg closest_so_far_outone_rsci_bcwt;
  input [46:0] closest_so_far_outone_rsci_idat;


  // Interconnect Declarations
  reg [46:0] closest_so_far_outone_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_outone_rsci_wen_comp = (~ closest_so_far_outone_rsci_oswt)
      | closest_so_far_outone_rsci_biwt | closest_so_far_outone_rsci_bcwt;
  assign closest_so_far_outone_rsci_idat_mxwt = MUX_v_47_2_2(closest_so_far_outone_rsci_idat,
      closest_so_far_outone_rsci_idat_bfwt, closest_so_far_outone_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_outone_rsci_bcwt <= 1'b0;
    end
    else begin
      closest_so_far_outone_rsci_bcwt <= ~((~(closest_so_far_outone_rsci_bcwt | closest_so_far_outone_rsci_biwt))
          | closest_so_far_outone_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_outone_rsci_idat_bfwt <= 47'b00000000000000000000000000000000000000000000000;
    end
    else if ( ~ closest_so_far_outone_rsci_bcwt ) begin
      closest_so_far_outone_rsci_idat_bfwt <= closest_so_far_outone_rsci_idat_mxwt;
    end
  end

  function automatic [46:0] MUX_v_47_2_2;
    input [46:0] input_0;
    input [46:0] input_1;
    input [0:0] sel;
    reg [46:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_47_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_ctrl (
  hit_wen, closest_so_far_outone_rsci_oswt, closest_so_far_outone_rsci_biwt, closest_so_far_outone_rsci_bdwt,
      closest_so_far_outone_rsci_bcwt, closest_so_far_outone_rsci_irdy_hit_sct, closest_so_far_outone_rsci_ivld
);
  input hit_wen;
  input closest_so_far_outone_rsci_oswt;
  output closest_so_far_outone_rsci_biwt;
  output closest_so_far_outone_rsci_bdwt;
  input closest_so_far_outone_rsci_bcwt;
  output closest_so_far_outone_rsci_irdy_hit_sct;
  input closest_so_far_outone_rsci_ivld;


  // Interconnect Declarations
  wire closest_so_far_outone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign closest_so_far_outone_rsci_bdwt = closest_so_far_outone_rsci_oswt & hit_wen;
  assign closest_so_far_outone_rsci_biwt = closest_so_far_outone_rsci_ogwt & closest_so_far_outone_rsci_ivld;
  assign closest_so_far_outone_rsci_ogwt = closest_so_far_outone_rsci_oswt & (~ closest_so_far_outone_rsci_bcwt);
  assign closest_so_far_outone_rsci_irdy_hit_sct = closest_so_far_outone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_dp (
  clk, arst_n, rec_quad_outtwo_rsci_oswt, rec_quad_outtwo_rsci_wen_comp, rec_quad_outtwo_rsci_idat_mxwt,
      rec_quad_outtwo_rsci_biwt, rec_quad_outtwo_rsci_bdwt, rec_quad_outtwo_rsci_bcwt,
      rec_quad_outtwo_rsci_idat
);
  input clk;
  input arst_n;
  input rec_quad_outtwo_rsci_oswt;
  output rec_quad_outtwo_rsci_wen_comp;
  output [225:0] rec_quad_outtwo_rsci_idat_mxwt;
  input rec_quad_outtwo_rsci_biwt;
  input rec_quad_outtwo_rsci_bdwt;
  output rec_quad_outtwo_rsci_bcwt;
  reg rec_quad_outtwo_rsci_bcwt;
  input [225:0] rec_quad_outtwo_rsci_idat;


  // Interconnect Declarations
  reg [225:0] rec_quad_outtwo_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_outtwo_rsci_wen_comp = (~ rec_quad_outtwo_rsci_oswt) | rec_quad_outtwo_rsci_biwt
      | rec_quad_outtwo_rsci_bcwt;
  assign rec_quad_outtwo_rsci_idat_mxwt = MUX_v_226_2_2(rec_quad_outtwo_rsci_idat,
      rec_quad_outtwo_rsci_idat_bfwt, rec_quad_outtwo_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_outtwo_rsci_bcwt <= 1'b0;
    end
    else begin
      rec_quad_outtwo_rsci_bcwt <= ~((~(rec_quad_outtwo_rsci_bcwt | rec_quad_outtwo_rsci_biwt))
          | rec_quad_outtwo_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_outtwo_rsci_idat_bfwt <= 226'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ rec_quad_outtwo_rsci_bcwt ) begin
      rec_quad_outtwo_rsci_idat_bfwt <= rec_quad_outtwo_rsci_idat_mxwt;
    end
  end

  function automatic [225:0] MUX_v_226_2_2;
    input [225:0] input_0;
    input [225:0] input_1;
    input [0:0] sel;
    reg [225:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_226_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_ctrl (
  hit_wen, rec_quad_outtwo_rsci_oswt, rec_quad_outtwo_rsci_biwt, rec_quad_outtwo_rsci_bdwt,
      rec_quad_outtwo_rsci_bcwt, rec_quad_outtwo_rsci_irdy_hit_sct, rec_quad_outtwo_rsci_ivld
);
  input hit_wen;
  input rec_quad_outtwo_rsci_oswt;
  output rec_quad_outtwo_rsci_biwt;
  output rec_quad_outtwo_rsci_bdwt;
  input rec_quad_outtwo_rsci_bcwt;
  output rec_quad_outtwo_rsci_irdy_hit_sct;
  input rec_quad_outtwo_rsci_ivld;


  // Interconnect Declarations
  wire rec_quad_outtwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_outtwo_rsci_bdwt = rec_quad_outtwo_rsci_oswt & hit_wen;
  assign rec_quad_outtwo_rsci_biwt = rec_quad_outtwo_rsci_ogwt & rec_quad_outtwo_rsci_ivld;
  assign rec_quad_outtwo_rsci_ogwt = rec_quad_outtwo_rsci_oswt & (~ rec_quad_outtwo_rsci_bcwt);
  assign rec_quad_outtwo_rsci_irdy_hit_sct = rec_quad_outtwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_dp (
  clk, arst_n, rec_quad_outone_rsci_oswt, rec_quad_outone_rsci_wen_comp, rec_quad_outone_rsci_idat_mxwt,
      rec_quad_outone_rsci_biwt, rec_quad_outone_rsci_bdwt, rec_quad_outone_rsci_bcwt,
      rec_quad_outone_rsci_idat
);
  input clk;
  input arst_n;
  input rec_quad_outone_rsci_oswt;
  output rec_quad_outone_rsci_wen_comp;
  output [225:0] rec_quad_outone_rsci_idat_mxwt;
  input rec_quad_outone_rsci_biwt;
  input rec_quad_outone_rsci_bdwt;
  output rec_quad_outone_rsci_bcwt;
  reg rec_quad_outone_rsci_bcwt;
  input [225:0] rec_quad_outone_rsci_idat;


  // Interconnect Declarations
  reg [225:0] rec_quad_outone_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_outone_rsci_wen_comp = (~ rec_quad_outone_rsci_oswt) | rec_quad_outone_rsci_biwt
      | rec_quad_outone_rsci_bcwt;
  assign rec_quad_outone_rsci_idat_mxwt = MUX_v_226_2_2(rec_quad_outone_rsci_idat,
      rec_quad_outone_rsci_idat_bfwt, rec_quad_outone_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_outone_rsci_bcwt <= 1'b0;
    end
    else begin
      rec_quad_outone_rsci_bcwt <= ~((~(rec_quad_outone_rsci_bcwt | rec_quad_outone_rsci_biwt))
          | rec_quad_outone_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_outone_rsci_idat_bfwt <= 226'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ rec_quad_outone_rsci_bcwt ) begin
      rec_quad_outone_rsci_idat_bfwt <= rec_quad_outone_rsci_idat_mxwt;
    end
  end

  function automatic [225:0] MUX_v_226_2_2;
    input [225:0] input_0;
    input [225:0] input_1;
    input [0:0] sel;
    reg [225:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_226_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_ctrl (
  hit_wen, rec_quad_outone_rsci_oswt, rec_quad_outone_rsci_biwt, rec_quad_outone_rsci_bdwt,
      rec_quad_outone_rsci_bcwt, rec_quad_outone_rsci_irdy_hit_sct, rec_quad_outone_rsci_ivld
);
  input hit_wen;
  input rec_quad_outone_rsci_oswt;
  output rec_quad_outone_rsci_biwt;
  output rec_quad_outone_rsci_bdwt;
  input rec_quad_outone_rsci_bcwt;
  output rec_quad_outone_rsci_irdy_hit_sct;
  input rec_quad_outone_rsci_ivld;


  // Interconnect Declarations
  wire rec_quad_outone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rec_quad_outone_rsci_bdwt = rec_quad_outone_rsci_oswt & hit_wen;
  assign rec_quad_outone_rsci_biwt = rec_quad_outone_rsci_ogwt & rec_quad_outone_rsci_ivld;
  assign rec_quad_outone_rsci_ogwt = rec_quad_outone_rsci_oswt & (~ rec_quad_outone_rsci_bcwt);
  assign rec_quad_outone_rsci_irdy_hit_sct = rec_quad_outone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_dp
    (
  clk, arst_n, quad_hit_anything_outtwo_rsci_oswt, quad_hit_anything_outtwo_rsci_wen_comp,
      quad_hit_anything_outtwo_rsci_idat_mxwt, quad_hit_anything_outtwo_rsci_biwt,
      quad_hit_anything_outtwo_rsci_bdwt, quad_hit_anything_outtwo_rsci_bcwt, quad_hit_anything_outtwo_rsci_idat
);
  input clk;
  input arst_n;
  input quad_hit_anything_outtwo_rsci_oswt;
  output quad_hit_anything_outtwo_rsci_wen_comp;
  output quad_hit_anything_outtwo_rsci_idat_mxwt;
  input quad_hit_anything_outtwo_rsci_biwt;
  input quad_hit_anything_outtwo_rsci_bdwt;
  output quad_hit_anything_outtwo_rsci_bcwt;
  reg quad_hit_anything_outtwo_rsci_bcwt;
  input quad_hit_anything_outtwo_rsci_idat;


  // Interconnect Declarations
  reg quad_hit_anything_outtwo_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_outtwo_rsci_wen_comp = (~ quad_hit_anything_outtwo_rsci_oswt)
      | quad_hit_anything_outtwo_rsci_biwt | quad_hit_anything_outtwo_rsci_bcwt;
  assign quad_hit_anything_outtwo_rsci_idat_mxwt = MUX_s_1_2_2(quad_hit_anything_outtwo_rsci_idat,
      quad_hit_anything_outtwo_rsci_idat_bfwt, quad_hit_anything_outtwo_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_outtwo_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_hit_anything_outtwo_rsci_bcwt <= ~((~(quad_hit_anything_outtwo_rsci_bcwt
          | quad_hit_anything_outtwo_rsci_biwt)) | quad_hit_anything_outtwo_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_outtwo_rsci_idat_bfwt <= 1'b0;
    end
    else if ( ~ quad_hit_anything_outtwo_rsci_bcwt ) begin
      quad_hit_anything_outtwo_rsci_idat_bfwt <= quad_hit_anything_outtwo_rsci_idat_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_ctrl
    (
  hit_wen, quad_hit_anything_outtwo_rsci_oswt, quad_hit_anything_outtwo_rsci_biwt,
      quad_hit_anything_outtwo_rsci_bdwt, quad_hit_anything_outtwo_rsci_bcwt, quad_hit_anything_outtwo_rsci_irdy_hit_sct,
      quad_hit_anything_outtwo_rsci_ivld
);
  input hit_wen;
  input quad_hit_anything_outtwo_rsci_oswt;
  output quad_hit_anything_outtwo_rsci_biwt;
  output quad_hit_anything_outtwo_rsci_bdwt;
  input quad_hit_anything_outtwo_rsci_bcwt;
  output quad_hit_anything_outtwo_rsci_irdy_hit_sct;
  input quad_hit_anything_outtwo_rsci_ivld;


  // Interconnect Declarations
  wire quad_hit_anything_outtwo_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_outtwo_rsci_bdwt = quad_hit_anything_outtwo_rsci_oswt
      & hit_wen;
  assign quad_hit_anything_outtwo_rsci_biwt = quad_hit_anything_outtwo_rsci_ogwt
      & quad_hit_anything_outtwo_rsci_ivld;
  assign quad_hit_anything_outtwo_rsci_ogwt = quad_hit_anything_outtwo_rsci_oswt
      & (~ quad_hit_anything_outtwo_rsci_bcwt);
  assign quad_hit_anything_outtwo_rsci_irdy_hit_sct = quad_hit_anything_outtwo_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_dp
    (
  clk, arst_n, quad_hit_anything_outone_rsci_oswt, quad_hit_anything_outone_rsci_wen_comp,
      quad_hit_anything_outone_rsci_idat_mxwt, quad_hit_anything_outone_rsci_biwt,
      quad_hit_anything_outone_rsci_bdwt, quad_hit_anything_outone_rsci_bcwt, quad_hit_anything_outone_rsci_idat
);
  input clk;
  input arst_n;
  input quad_hit_anything_outone_rsci_oswt;
  output quad_hit_anything_outone_rsci_wen_comp;
  output quad_hit_anything_outone_rsci_idat_mxwt;
  input quad_hit_anything_outone_rsci_biwt;
  input quad_hit_anything_outone_rsci_bdwt;
  output quad_hit_anything_outone_rsci_bcwt;
  reg quad_hit_anything_outone_rsci_bcwt;
  input quad_hit_anything_outone_rsci_idat;


  // Interconnect Declarations
  reg quad_hit_anything_outone_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_outone_rsci_wen_comp = (~ quad_hit_anything_outone_rsci_oswt)
      | quad_hit_anything_outone_rsci_biwt | quad_hit_anything_outone_rsci_bcwt;
  assign quad_hit_anything_outone_rsci_idat_mxwt = MUX_s_1_2_2(quad_hit_anything_outone_rsci_idat,
      quad_hit_anything_outone_rsci_idat_bfwt, quad_hit_anything_outone_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_outone_rsci_bcwt <= 1'b0;
    end
    else begin
      quad_hit_anything_outone_rsci_bcwt <= ~((~(quad_hit_anything_outone_rsci_bcwt
          | quad_hit_anything_outone_rsci_biwt)) | quad_hit_anything_outone_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_outone_rsci_idat_bfwt <= 1'b0;
    end
    else if ( ~ quad_hit_anything_outone_rsci_bcwt ) begin
      quad_hit_anything_outone_rsci_idat_bfwt <= quad_hit_anything_outone_rsci_idat_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_ctrl
    (
  hit_wen, quad_hit_anything_outone_rsci_oswt, quad_hit_anything_outone_rsci_biwt,
      quad_hit_anything_outone_rsci_bdwt, quad_hit_anything_outone_rsci_bcwt, quad_hit_anything_outone_rsci_irdy_hit_sct,
      quad_hit_anything_outone_rsci_ivld
);
  input hit_wen;
  input quad_hit_anything_outone_rsci_oswt;
  output quad_hit_anything_outone_rsci_biwt;
  output quad_hit_anything_outone_rsci_bdwt;
  input quad_hit_anything_outone_rsci_bcwt;
  output quad_hit_anything_outone_rsci_irdy_hit_sct;
  input quad_hit_anything_outone_rsci_ivld;


  // Interconnect Declarations
  wire quad_hit_anything_outone_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign quad_hit_anything_outone_rsci_bdwt = quad_hit_anything_outone_rsci_oswt
      & hit_wen;
  assign quad_hit_anything_outone_rsci_biwt = quad_hit_anything_outone_rsci_ogwt
      & quad_hit_anything_outone_rsci_ivld;
  assign quad_hit_anything_outone_rsci_ogwt = quad_hit_anything_outone_rsci_oswt
      & (~ quad_hit_anything_outone_rsci_bcwt);
  assign quad_hit_anything_outone_rsci_irdy_hit_sct = quad_hit_anything_outone_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
    (
  clk, arst_n, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_idat_mxwt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  input accumalated_color_chan_in_rsci_biwt;
  input accumalated_color_chan_in_rsci_bdwt;
  output accumalated_color_chan_in_rsci_bcwt;
  reg accumalated_color_chan_in_rsci_bcwt;
  input [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] accumalated_color_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_wen_comp = (~ accumalated_color_chan_in_rsci_oswt)
      | accumalated_color_chan_in_rsci_biwt | accumalated_color_chan_in_rsci_bcwt;
  assign accumalated_color_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(accumalated_color_chan_in_rsci_idat,
      accumalated_color_chan_in_rsci_idat_bfwt, accumalated_color_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_chan_in_rsci_bcwt <= ~((~(accumalated_color_chan_in_rsci_bcwt
          | accumalated_color_chan_in_rsci_biwt)) | accumalated_color_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ accumalated_color_chan_in_rsci_bcwt ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
    (
  hit_wen, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_irdy_hit_sct,
      accumalated_color_chan_in_rsci_ivld
);
  input hit_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_biwt;
  output accumalated_color_chan_in_rsci_bdwt;
  input accumalated_color_chan_in_rsci_bcwt;
  output accumalated_color_chan_in_rsci_irdy_hit_sct;
  input accumalated_color_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_bdwt = accumalated_color_chan_in_rsci_oswt
      & hit_wen;
  assign accumalated_color_chan_in_rsci_biwt = accumalated_color_chan_in_rsci_ogwt
      & accumalated_color_chan_in_rsci_ivld;
  assign accumalated_color_chan_in_rsci_ogwt = accumalated_color_chan_in_rsci_oswt
      & (~ accumalated_color_chan_in_rsci_bcwt);
  assign accumalated_color_chan_in_rsci_irdy_hit_sct = accumalated_color_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp (
  clk, arst_n, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;
  input attenuation_chan_in_rsci_biwt;
  input attenuation_chan_in_rsci_bdwt;
  output attenuation_chan_in_rsci_bcwt;
  reg attenuation_chan_in_rsci_bcwt;
  input [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] attenuation_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_wen_comp = (~ attenuation_chan_in_rsci_oswt) |
      attenuation_chan_in_rsci_biwt | attenuation_chan_in_rsci_bcwt;
  assign attenuation_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(attenuation_chan_in_rsci_idat,
      attenuation_chan_in_rsci_idat_bfwt, attenuation_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_in_rsci_bcwt <= ~((~(attenuation_chan_in_rsci_bcwt | attenuation_chan_in_rsci_biwt))
          | attenuation_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ attenuation_chan_in_rsci_bcwt ) begin
      attenuation_chan_in_rsci_idat_bfwt <= attenuation_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl (
  hit_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_irdy_hit_sct, attenuation_chan_in_rsci_ivld
);
  input hit_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_biwt;
  output attenuation_chan_in_rsci_bdwt;
  input attenuation_chan_in_rsci_bcwt;
  output attenuation_chan_in_rsci_irdy_hit_sct;
  input attenuation_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_bdwt = attenuation_chan_in_rsci_oswt & hit_wen;
  assign attenuation_chan_in_rsci_biwt = attenuation_chan_in_rsci_ogwt & attenuation_chan_in_rsci_ivld;
  assign attenuation_chan_in_rsci_ogwt = attenuation_chan_in_rsci_oswt & (~ attenuation_chan_in_rsci_bcwt);
  assign attenuation_chan_in_rsci_irdy_hit_sct = attenuation_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_params_in_rsci_params_in_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_params_in_rsci_params_in_wait_dp (
  clk, arst_n, params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt,
      params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt, params_in_rsci_idat
);
  input clk;
  input arst_n;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [80:0] params_in_rsci_idat_mxwt;
  input params_in_rsci_biwt;
  input params_in_rsci_bdwt;
  output params_in_rsci_bcwt;
  reg params_in_rsci_bcwt;
  input [92:0] params_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] params_in_rsci_idat_bfwt_91_11;
  wire [80:0] params_in_rsci_idat_mxwt_opt_91_11;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_wen_comp = (~ params_in_rsci_oswt) | params_in_rsci_biwt
      | params_in_rsci_bcwt;
  assign params_in_rsci_idat_mxwt_opt_91_11 = MUX_v_81_2_2((params_in_rsci_idat[91:11]),
      params_in_rsci_idat_bfwt_91_11, params_in_rsci_bcwt);
  assign params_in_rsci_idat_mxwt = params_in_rsci_idat_mxwt_opt_91_11;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_bcwt <= 1'b0;
    end
    else begin
      params_in_rsci_bcwt <= ~((~(params_in_rsci_bcwt | params_in_rsci_biwt)) | params_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_idat_bfwt_91_11 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ params_in_rsci_bcwt ) begin
      params_in_rsci_idat_bfwt_91_11 <= params_in_rsci_idat_mxwt_opt_91_11;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_params_in_rsci_params_in_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_params_in_rsci_params_in_wait_ctrl (
  hit_wen, params_in_rsci_oswt, params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt,
      params_in_rsci_irdy_hit_sct, params_in_rsci_ivld
);
  input hit_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_biwt;
  output params_in_rsci_bdwt;
  input params_in_rsci_bcwt;
  output params_in_rsci_irdy_hit_sct;
  input params_in_rsci_ivld;


  // Interconnect Declarations
  wire params_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_bdwt = params_in_rsci_oswt & hit_wen;
  assign params_in_rsci_biwt = params_in_rsci_ogwt & params_in_rsci_ivld;
  assign params_in_rsci_ogwt = params_in_rsci_oswt & (~ params_in_rsci_bcwt);
  assign params_in_rsci_irdy_hit_sct = params_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_in_rsci_ray_in_wait_dp
// ------------------------------------------------------------------


module WorldHit_hit_ray_in_rsci_ray_in_wait_dp (
  clk, arst_n, ray_in_rsci_oswt, ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt, ray_in_rsci_biwt,
      ray_in_rsci_bdwt, ray_in_rsci_bcwt, ray_in_rsci_idat
);
  input clk;
  input arst_n;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [164:0] ray_in_rsci_idat_mxwt;
  input ray_in_rsci_biwt;
  input ray_in_rsci_bdwt;
  output ray_in_rsci_bcwt;
  reg ray_in_rsci_bcwt;
  input [165:0] ray_in_rsci_idat;


  // Interconnect Declarations
  reg [164:0] ray_in_rsci_idat_bfwt_164_0;
  wire [164:0] ray_in_rsci_idat_mxwt_opt_164_0;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_wen_comp = (~ ray_in_rsci_oswt) | ray_in_rsci_biwt | ray_in_rsci_bcwt;
  assign ray_in_rsci_idat_mxwt_opt_164_0 = MUX_v_165_2_2((ray_in_rsci_idat[164:0]),
      ray_in_rsci_idat_bfwt_164_0, ray_in_rsci_bcwt);
  assign ray_in_rsci_idat_mxwt = ray_in_rsci_idat_mxwt_opt_164_0;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_in_rsci_bcwt <= ~((~(ray_in_rsci_bcwt | ray_in_rsci_biwt)) | ray_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_idat_bfwt_164_0 <= 165'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_in_rsci_bcwt ) begin
      ray_in_rsci_idat_bfwt_164_0 <= ray_in_rsci_idat_mxwt_opt_164_0;
    end
  end

  function automatic [164:0] MUX_v_165_2_2;
    input [164:0] input_0;
    input [164:0] input_1;
    input [0:0] sel;
    reg [164:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_165_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_in_rsci_ray_in_wait_ctrl
// ------------------------------------------------------------------


module WorldHit_hit_ray_in_rsci_ray_in_wait_ctrl (
  hit_wen, ray_in_rsci_oswt, ray_in_rsci_biwt, ray_in_rsci_bdwt, ray_in_rsci_bcwt,
      ray_in_rsci_irdy_hit_sct, ray_in_rsci_ivld
);
  input hit_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_biwt;
  output ray_in_rsci_bdwt;
  input ray_in_rsci_bcwt;
  output ray_in_rsci_irdy_hit_sct;
  input ray_in_rsci_ivld;


  // Interconnect Declarations
  wire ray_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_bdwt = ray_in_rsci_oswt & hit_wen;
  assign ray_in_rsci_biwt = ray_in_rsci_ogwt & ray_in_rsci_ivld;
  assign ray_in_rsci_ogwt = ray_in_rsci_oswt & (~ ray_in_rsci_bcwt);
  assign ray_in_rsci_irdy_hit_sct = ray_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_scatter_fsm
//  FSM Module
// ------------------------------------------------------------------


module MaterialScatter_scatter_scatter_fsm (
  clk, arst_n, scatter_wen, fsm_output, main_C_4_tr0, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0,
      main_C_7_tr0, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1_tr0
);
  input clk;
  input arst_n;
  input scatter_wen;
  output [20:0] fsm_output;
  reg [20:0] fsm_output;
  input main_C_4_tr0;
  input ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0;
  input main_C_7_tr0;
  input ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1_tr0;


  // FSM State Type Declaration for MaterialScatter_scatter_scatter_fsm_1
  parameter
    scatter_rlp_C_0 = 5'd0,
    main_C_0 = 5'd1,
    main_C_1 = 5'd2,
    main_C_2 = 5'd3,
    main_C_3 = 5'd4,
    main_C_4 = 5'd5,
    ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0 = 5'd6,
    ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1 = 5'd7,
    ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2 = 5'd8,
    main_C_5 = 5'd9,
    main_C_6 = 5'd10,
    main_C_7 = 5'd11,
    ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0 = 5'd12,
    ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1 = 5'd13,
    main_C_8 = 5'd14,
    main_C_9 = 5'd15,
    main_C_10 = 5'd16,
    main_C_11 = 5'd17,
    main_C_12 = 5'd18,
    main_C_13 = 5'd19,
    main_C_14 = 5'd20;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : MaterialScatter_scatter_scatter_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 21'b000000000000000000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 21'b000000000000000000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 21'b000000000000000001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 21'b000000000000000010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 21'b000000000000000100000;
        if ( main_C_4_tr0 ) begin
          state_var_NS = main_C_5;
        end
        else begin
          state_var_NS = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0;
        end
      end
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0 :
          begin
        fsm_output = 21'b000000000000001000000;
        state_var_NS = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1;
      end
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1 :
          begin
        fsm_output = 21'b000000000000010000000;
        state_var_NS = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2;
      end
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2 :
          begin
        fsm_output = 21'b000000000000100000000;
        if ( ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0
            ) begin
          state_var_NS = main_C_5;
        end
        else begin
          state_var_NS = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0;
        end
      end
      main_C_5 : begin
        fsm_output = 21'b000000000001000000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 21'b000000000010000000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 21'b000000000100000000000;
        if ( main_C_7_tr0 ) begin
          state_var_NS = main_C_8;
        end
        else begin
          state_var_NS = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0;
        end
      end
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0 :
          begin
        fsm_output = 21'b000000001000000000000;
        state_var_NS = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1;
      end
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1 :
          begin
        fsm_output = 21'b000000010000000000000;
        if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1_tr0
            ) begin
          state_var_NS = main_C_8;
        end
        else begin
          state_var_NS = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_0;
        end
      end
      main_C_8 : begin
        fsm_output = 21'b000000100000000000000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 21'b000001000000000000000;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 21'b000010000000000000000;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 21'b000100000000000000000;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 21'b001000000000000000000;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 21'b010000000000000000000;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 21'b100000000000000000000;
        state_var_NS = main_C_0;
      end
      // scatter_rlp_C_0
      default : begin
        fsm_output = 21'b000000000000000000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= scatter_rlp_C_0;
    end
    else if ( scatter_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_staller
// ------------------------------------------------------------------


module MaterialScatter_scatter_staller (
  scatter_wen, ray_in_rsci_wen_comp, hit_in_rsci_wen_comp, attenuation_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_wen_comp, isHit_rsci_wen_comp, attenuation_chan_out_rsci_wen_comp,
      accumalated_color_out_rsci_wen_comp, ray_out_rsci_wen_comp
);
  output scatter_wen;
  input ray_in_rsci_wen_comp;
  input hit_in_rsci_wen_comp;
  input attenuation_chan_in_rsci_wen_comp;
  input accumalated_color_chan_in_rsci_wen_comp;
  input isHit_rsci_wen_comp;
  input attenuation_chan_out_rsci_wen_comp;
  input accumalated_color_out_rsci_wen_comp;
  input ray_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign scatter_wen = ray_in_rsci_wen_comp & hit_in_rsci_wen_comp & attenuation_chan_in_rsci_wen_comp
      & accumalated_color_chan_in_rsci_wen_comp & isHit_rsci_wen_comp & attenuation_chan_out_rsci_wen_comp
      & accumalated_color_out_rsci_wen_comp & ray_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_wait_dp (
  clk, arst_n, ensig_cgo_iro, lambertianScatter_rand_unit_run_xs_mul_cmp_en, lambertianScatter_rand_unit_run_xs_mul_cmp_z,
      else_if_mul_cmp_z, scatter_wen, ensig_cgo, lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg,
      else_if_mul_cmp_z_oreg
);
  input clk;
  input arst_n;
  input ensig_cgo_iro;
  output lambertianScatter_rand_unit_run_xs_mul_cmp_en;
  input [65:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z;
  input [48:0] else_if_mul_cmp_z;
  input scatter_wen;
  input ensig_cgo;
  output [33:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg;
  output [26:0] else_if_mul_cmp_z_oreg;


  // Interconnect Declarations
  reg [33:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg_pconst_65_32;
  reg [26:0] else_if_mul_cmp_z_oreg_pconst_48_22;


  // Interconnect Declarations for Component Instantiations 
  assign lambertianScatter_rand_unit_run_xs_mul_cmp_en = ~(scatter_wen & (ensig_cgo
      | ensig_cgo_iro));
  assign lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg = lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg_pconst_65_32;
  assign else_if_mul_cmp_z_oreg = else_if_mul_cmp_z_oreg_pconst_48_22;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg_pconst_65_32 <= 34'b0000000000000000000000000000000000;
    end
    else if ( ~ lambertianScatter_rand_unit_run_xs_mul_cmp_en ) begin
      lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg_pconst_65_32 <= lambertianScatter_rand_unit_run_xs_mul_cmp_z[65:32];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      else_if_mul_cmp_z_oreg_pconst_48_22 <= 27'b000000000000000000000000000;
    end
    else if ( scatter_wen ) begin
      else_if_mul_cmp_z_oreg_pconst_48_22 <= else_if_mul_cmp_z[48:22];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_out_rsci_ray_out_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_out_rsci_ray_out_wait_dp (
  clk, arst_n, ray_out_rsci_oswt, ray_out_rsci_wen_comp, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input ray_out_rsci_biwt;
  input ray_out_rsci_bdwt;
  output ray_out_rsci_bcwt;
  reg ray_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_wen_comp = (~ ray_out_rsci_oswt) | ray_out_rsci_biwt | ray_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_rsci_bcwt <= ~((~(ray_out_rsci_bcwt | ray_out_rsci_biwt)) | ray_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_out_rsci_ray_out_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_out_rsci_ray_out_wait_ctrl (
  scatter_wen, ray_out_rsci_oswt, ray_out_rsci_irdy, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt, ray_out_rsci_ivld_scatter_sct
);
  input scatter_wen;
  input ray_out_rsci_oswt;
  input ray_out_rsci_irdy;
  output ray_out_rsci_biwt;
  output ray_out_rsci_bdwt;
  input ray_out_rsci_bcwt;
  output ray_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations
  wire ray_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_bdwt = ray_out_rsci_oswt & scatter_wen;
  assign ray_out_rsci_biwt = ray_out_rsci_ogwt & ray_out_rsci_irdy;
  assign ray_out_rsci_ogwt = ray_out_rsci_oswt & (~ ray_out_rsci_bcwt);
  assign ray_out_rsci_ivld_scatter_sct = ray_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_dp
    (
  clk, arst_n, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_biwt, accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input accumalated_color_out_rsci_biwt;
  input accumalated_color_out_rsci_bdwt;
  output accumalated_color_out_rsci_bcwt;
  reg accumalated_color_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_wen_comp = (~ accumalated_color_out_rsci_oswt)
      | accumalated_color_out_rsci_biwt | accumalated_color_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_out_rsci_bcwt <= ~((~(accumalated_color_out_rsci_bcwt | accumalated_color_out_rsci_biwt))
          | accumalated_color_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
    (
  scatter_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_irdy,
      accumalated_color_out_rsci_biwt, accumalated_color_out_rsci_bdwt, accumalated_color_out_rsci_bcwt,
      accumalated_color_out_rsci_ivld_scatter_sct
);
  input scatter_wen;
  input accumalated_color_out_rsci_oswt;
  input accumalated_color_out_rsci_irdy;
  output accumalated_color_out_rsci_biwt;
  output accumalated_color_out_rsci_bdwt;
  input accumalated_color_out_rsci_bcwt;
  output accumalated_color_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_out_rsci_bdwt = accumalated_color_out_rsci_oswt & scatter_wen;
  assign accumalated_color_out_rsci_biwt = accumalated_color_out_rsci_ogwt & accumalated_color_out_rsci_irdy;
  assign accumalated_color_out_rsci_ogwt = accumalated_color_out_rsci_oswt & (~ accumalated_color_out_rsci_bcwt);
  assign accumalated_color_out_rsci_ivld_scatter_sct = accumalated_color_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp
    (
  clk, arst_n, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_biwt, attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input attenuation_chan_out_rsci_biwt;
  input attenuation_chan_out_rsci_bdwt;
  output attenuation_chan_out_rsci_bcwt;
  reg attenuation_chan_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_wen_comp = (~ attenuation_chan_out_rsci_oswt)
      | attenuation_chan_out_rsci_biwt | attenuation_chan_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_out_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_out_rsci_bcwt <= ~((~(attenuation_chan_out_rsci_bcwt | attenuation_chan_out_rsci_biwt))
          | attenuation_chan_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl
    (
  scatter_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_irdy, attenuation_chan_out_rsci_biwt,
      attenuation_chan_out_rsci_bdwt, attenuation_chan_out_rsci_bcwt, attenuation_chan_out_rsci_ivld_scatter_sct
);
  input scatter_wen;
  input attenuation_chan_out_rsci_oswt;
  input attenuation_chan_out_rsci_irdy;
  output attenuation_chan_out_rsci_biwt;
  output attenuation_chan_out_rsci_bdwt;
  input attenuation_chan_out_rsci_bcwt;
  output attenuation_chan_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_out_rsci_bdwt = attenuation_chan_out_rsci_oswt & scatter_wen;
  assign attenuation_chan_out_rsci_biwt = attenuation_chan_out_rsci_ogwt & attenuation_chan_out_rsci_irdy;
  assign attenuation_chan_out_rsci_ogwt = attenuation_chan_out_rsci_oswt & (~ attenuation_chan_out_rsci_bcwt);
  assign attenuation_chan_out_rsci_ivld_scatter_sct = attenuation_chan_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_isHit_rsci_isHit_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_isHit_rsci_isHit_wait_dp (
  clk, arst_n, isHit_rsci_oswt, isHit_rsci_wen_comp, isHit_rsci_idat_mxwt, isHit_rsci_biwt,
      isHit_rsci_bdwt, isHit_rsci_bcwt, isHit_rsci_idat
);
  input clk;
  input arst_n;
  input isHit_rsci_oswt;
  output isHit_rsci_wen_comp;
  output isHit_rsci_idat_mxwt;
  input isHit_rsci_biwt;
  input isHit_rsci_bdwt;
  output isHit_rsci_bcwt;
  reg isHit_rsci_bcwt;
  input isHit_rsci_idat;


  // Interconnect Declarations
  reg isHit_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign isHit_rsci_wen_comp = (~ isHit_rsci_oswt) | isHit_rsci_biwt | isHit_rsci_bcwt;
  assign isHit_rsci_idat_mxwt = MUX_s_1_2_2(isHit_rsci_idat, isHit_rsci_idat_bfwt,
      isHit_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      isHit_rsci_bcwt <= 1'b0;
    end
    else begin
      isHit_rsci_bcwt <= ~((~(isHit_rsci_bcwt | isHit_rsci_biwt)) | isHit_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      isHit_rsci_idat_bfwt <= 1'b0;
    end
    else if ( ~ isHit_rsci_bcwt ) begin
      isHit_rsci_idat_bfwt <= isHit_rsci_idat_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_isHit_rsci_isHit_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_isHit_rsci_isHit_wait_ctrl (
  scatter_wen, isHit_rsci_oswt, isHit_rsci_biwt, isHit_rsci_bdwt, isHit_rsci_bcwt,
      isHit_rsci_irdy_scatter_sct, isHit_rsci_ivld
);
  input scatter_wen;
  input isHit_rsci_oswt;
  output isHit_rsci_biwt;
  output isHit_rsci_bdwt;
  input isHit_rsci_bcwt;
  output isHit_rsci_irdy_scatter_sct;
  input isHit_rsci_ivld;


  // Interconnect Declarations
  wire isHit_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign isHit_rsci_bdwt = isHit_rsci_oswt & scatter_wen;
  assign isHit_rsci_biwt = isHit_rsci_ogwt & isHit_rsci_ivld;
  assign isHit_rsci_ogwt = isHit_rsci_oswt & (~ isHit_rsci_bcwt);
  assign isHit_rsci_irdy_scatter_sct = isHit_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
    (
  clk, arst_n, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_wen_comp,
      accumalated_color_chan_in_rsci_idat_mxwt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  input accumalated_color_chan_in_rsci_biwt;
  input accumalated_color_chan_in_rsci_bdwt;
  output accumalated_color_chan_in_rsci_bcwt;
  reg accumalated_color_chan_in_rsci_bcwt;
  input [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] accumalated_color_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_wen_comp = (~ accumalated_color_chan_in_rsci_oswt)
      | accumalated_color_chan_in_rsci_biwt | accumalated_color_chan_in_rsci_bcwt;
  assign accumalated_color_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(accumalated_color_chan_in_rsci_idat,
      accumalated_color_chan_in_rsci_idat_bfwt, accumalated_color_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      accumalated_color_chan_in_rsci_bcwt <= ~((~(accumalated_color_chan_in_rsci_bcwt
          | accumalated_color_chan_in_rsci_biwt)) | accumalated_color_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ accumalated_color_chan_in_rsci_bcwt ) begin
      accumalated_color_chan_in_rsci_idat_bfwt <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
    (
  scatter_wen, accumalated_color_chan_in_rsci_oswt, accumalated_color_chan_in_rsci_biwt,
      accumalated_color_chan_in_rsci_bdwt, accumalated_color_chan_in_rsci_bcwt, accumalated_color_chan_in_rsci_irdy_scatter_sct,
      accumalated_color_chan_in_rsci_ivld
);
  input scatter_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_biwt;
  output accumalated_color_chan_in_rsci_bdwt;
  input accumalated_color_chan_in_rsci_bcwt;
  output accumalated_color_chan_in_rsci_irdy_scatter_sct;
  input accumalated_color_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumalated_color_chan_in_rsci_bdwt = accumalated_color_chan_in_rsci_oswt
      & scatter_wen;
  assign accumalated_color_chan_in_rsci_biwt = accumalated_color_chan_in_rsci_ogwt
      & accumalated_color_chan_in_rsci_ivld;
  assign accumalated_color_chan_in_rsci_ogwt = accumalated_color_chan_in_rsci_oswt
      & (~ accumalated_color_chan_in_rsci_bcwt);
  assign accumalated_color_chan_in_rsci_irdy_scatter_sct = accumalated_color_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp
    (
  clk, arst_n, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;
  input attenuation_chan_in_rsci_biwt;
  input attenuation_chan_in_rsci_bdwt;
  output attenuation_chan_in_rsci_bcwt;
  reg attenuation_chan_in_rsci_bcwt;
  input [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] attenuation_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_wen_comp = (~ attenuation_chan_in_rsci_oswt) |
      attenuation_chan_in_rsci_biwt | attenuation_chan_in_rsci_bcwt;
  assign attenuation_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(attenuation_chan_in_rsci_idat,
      attenuation_chan_in_rsci_idat_bfwt, attenuation_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      attenuation_chan_in_rsci_bcwt <= ~((~(attenuation_chan_in_rsci_bcwt | attenuation_chan_in_rsci_biwt))
          | attenuation_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ attenuation_chan_in_rsci_bcwt ) begin
      attenuation_chan_in_rsci_idat_bfwt <= attenuation_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl
    (
  scatter_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_biwt, attenuation_chan_in_rsci_bdwt,
      attenuation_chan_in_rsci_bcwt, attenuation_chan_in_rsci_irdy_scatter_sct, attenuation_chan_in_rsci_ivld
);
  input scatter_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_biwt;
  output attenuation_chan_in_rsci_bdwt;
  input attenuation_chan_in_rsci_bcwt;
  output attenuation_chan_in_rsci_irdy_scatter_sct;
  input attenuation_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign attenuation_chan_in_rsci_bdwt = attenuation_chan_in_rsci_oswt & scatter_wen;
  assign attenuation_chan_in_rsci_biwt = attenuation_chan_in_rsci_ogwt & attenuation_chan_in_rsci_ivld;
  assign attenuation_chan_in_rsci_ogwt = attenuation_chan_in_rsci_oswt & (~ attenuation_chan_in_rsci_bcwt);
  assign attenuation_chan_in_rsci_irdy_scatter_sct = attenuation_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_hit_in_rsci_hit_in_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_hit_in_rsci_hit_in_wait_dp (
  clk, arst_n, hit_in_rsci_oswt, hit_in_rsci_wen_comp, hit_in_rsci_idat_mxwt, hit_in_rsci_biwt,
      hit_in_rsci_bdwt, hit_in_rsci_bcwt, hit_in_rsci_idat
);
  input clk;
  input arst_n;
  input hit_in_rsci_oswt;
  output hit_in_rsci_wen_comp;
  output [225:0] hit_in_rsci_idat_mxwt;
  input hit_in_rsci_biwt;
  input hit_in_rsci_bdwt;
  output hit_in_rsci_bcwt;
  reg hit_in_rsci_bcwt;
  input [225:0] hit_in_rsci_idat;


  // Interconnect Declarations
  reg [225:0] hit_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign hit_in_rsci_wen_comp = (~ hit_in_rsci_oswt) | hit_in_rsci_biwt | hit_in_rsci_bcwt;
  assign hit_in_rsci_idat_mxwt = MUX_v_226_2_2(hit_in_rsci_idat, hit_in_rsci_idat_bfwt,
      hit_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      hit_in_rsci_bcwt <= 1'b0;
    end
    else begin
      hit_in_rsci_bcwt <= ~((~(hit_in_rsci_bcwt | hit_in_rsci_biwt)) | hit_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      hit_in_rsci_idat_bfwt <= 226'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ hit_in_rsci_bcwt ) begin
      hit_in_rsci_idat_bfwt <= hit_in_rsci_idat_mxwt;
    end
  end

  function automatic [225:0] MUX_v_226_2_2;
    input [225:0] input_0;
    input [225:0] input_1;
    input [0:0] sel;
    reg [225:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_226_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_hit_in_rsci_hit_in_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_hit_in_rsci_hit_in_wait_ctrl (
  scatter_wen, hit_in_rsci_oswt, hit_in_rsci_biwt, hit_in_rsci_bdwt, hit_in_rsci_bcwt,
      hit_in_rsci_irdy_scatter_sct, hit_in_rsci_ivld
);
  input scatter_wen;
  input hit_in_rsci_oswt;
  output hit_in_rsci_biwt;
  output hit_in_rsci_bdwt;
  input hit_in_rsci_bcwt;
  output hit_in_rsci_irdy_scatter_sct;
  input hit_in_rsci_ivld;


  // Interconnect Declarations
  wire hit_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign hit_in_rsci_bdwt = hit_in_rsci_oswt & scatter_wen;
  assign hit_in_rsci_biwt = hit_in_rsci_ogwt & hit_in_rsci_ivld;
  assign hit_in_rsci_ogwt = hit_in_rsci_oswt & (~ hit_in_rsci_bcwt);
  assign hit_in_rsci_irdy_scatter_sct = hit_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_in_rsci_ray_in_wait_dp
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_in_rsci_ray_in_wait_dp (
  clk, arst_n, ray_in_rsci_oswt, ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt, ray_in_rsci_biwt,
      ray_in_rsci_bdwt, ray_in_rsci_bcwt, ray_in_rsci_idat
);
  input clk;
  input arst_n;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [165:0] ray_in_rsci_idat_mxwt;
  input ray_in_rsci_biwt;
  input ray_in_rsci_bdwt;
  output ray_in_rsci_bcwt;
  reg ray_in_rsci_bcwt;
  input [165:0] ray_in_rsci_idat;


  // Interconnect Declarations
  reg [165:0] ray_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_wen_comp = (~ ray_in_rsci_oswt) | ray_in_rsci_biwt | ray_in_rsci_bcwt;
  assign ray_in_rsci_idat_mxwt = MUX_v_166_2_2(ray_in_rsci_idat, ray_in_rsci_idat_bfwt,
      ray_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_in_rsci_bcwt <= ~((~(ray_in_rsci_bcwt | ray_in_rsci_biwt)) | ray_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_in_rsci_bcwt ) begin
      ray_in_rsci_idat_bfwt <= ray_in_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_in_rsci_ray_in_wait_ctrl
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_in_rsci_ray_in_wait_ctrl (
  scatter_wen, ray_in_rsci_oswt, ray_in_rsci_biwt, ray_in_rsci_bdwt, ray_in_rsci_bcwt,
      ray_in_rsci_irdy_scatter_sct, ray_in_rsci_ivld
);
  input scatter_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_biwt;
  output ray_in_rsci_bdwt;
  input ray_in_rsci_bcwt;
  output ray_in_rsci_irdy_scatter_sct;
  input ray_in_rsci_ivld;


  // Interconnect Declarations
  wire ray_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_in_rsci_bdwt = ray_in_rsci_oswt & scatter_wen;
  assign ray_in_rsci_biwt = ray_in_rsci_ogwt & ray_in_rsci_ivld;
  assign ray_in_rsci_ogwt = ray_in_rsci_oswt & (~ ray_in_rsci_bcwt);
  assign ray_in_rsci_irdy_scatter_sct = ray_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ShaderFeedbackController_run_run_fsm (
  clk, arst_n, run_wen, fsm_output
);
  input clk;
  input arst_n;
  input run_wen;
  output [2:0] fsm_output;
  reg [2:0] fsm_output;


  // FSM State Type Declaration for ShaderFeedbackController_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    main_C_1 = 2'd2;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ShaderFeedbackController_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 3'b010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 3'b100;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 3'b001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_staller
// ------------------------------------------------------------------


module ShaderFeedbackController_run_staller (
  run_wen, ray_chan_in_rsci_wen_comp, ray_scattered_chan_rsci_wen_comp, params_in_rsci_wen_comp,
      color_chan_in_rsci_wen_comp, atten_chan_in_rsci_wen_comp, ray_out_rsci_wen_comp,
      params_out_rsci_wen_comp, color_chan_out_rsci_wen_comp, atten_chan_out_rsci_wen_comp,
      output_pxl_serial_rsci_wen_comp
);
  output run_wen;
  input ray_chan_in_rsci_wen_comp;
  input ray_scattered_chan_rsci_wen_comp;
  input params_in_rsci_wen_comp;
  input color_chan_in_rsci_wen_comp;
  input atten_chan_in_rsci_wen_comp;
  input ray_out_rsci_wen_comp;
  input params_out_rsci_wen_comp;
  input color_chan_out_rsci_wen_comp;
  input atten_chan_out_rsci_wen_comp;
  input output_pxl_serial_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = ray_chan_in_rsci_wen_comp & ray_scattered_chan_rsci_wen_comp &
      params_in_rsci_wen_comp & color_chan_in_rsci_wen_comp & atten_chan_in_rsci_wen_comp
      & ray_out_rsci_wen_comp & params_out_rsci_wen_comp & color_chan_out_rsci_wen_comp
      & atten_chan_out_rsci_wen_comp & output_pxl_serial_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp
    (
  clk, arst_n, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_wen_comp, output_pxl_serial_rsci_biwt,
      output_pxl_serial_rsci_bdwt, output_pxl_serial_rsci_bcwt
);
  input clk;
  input arst_n;
  input output_pxl_serial_rsci_oswt;
  output output_pxl_serial_rsci_wen_comp;
  input output_pxl_serial_rsci_biwt;
  input output_pxl_serial_rsci_bdwt;
  output output_pxl_serial_rsci_bcwt;
  reg output_pxl_serial_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_pxl_serial_rsci_wen_comp = (~ output_pxl_serial_rsci_oswt) | output_pxl_serial_rsci_biwt
      | output_pxl_serial_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_pxl_serial_rsci_bcwt <= 1'b0;
    end
    else begin
      output_pxl_serial_rsci_bcwt <= ~((~(output_pxl_serial_rsci_bcwt | output_pxl_serial_rsci_biwt))
          | output_pxl_serial_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl
    (
  run_wen, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_irdy, output_pxl_serial_rsci_biwt,
      output_pxl_serial_rsci_bdwt, output_pxl_serial_rsci_bcwt, output_pxl_serial_rsci_ivld_run_sct
);
  input run_wen;
  input output_pxl_serial_rsci_oswt;
  input output_pxl_serial_rsci_irdy;
  output output_pxl_serial_rsci_biwt;
  output output_pxl_serial_rsci_bdwt;
  input output_pxl_serial_rsci_bcwt;
  output output_pxl_serial_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire output_pxl_serial_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_pxl_serial_rsci_bdwt = output_pxl_serial_rsci_oswt & run_wen;
  assign output_pxl_serial_rsci_biwt = output_pxl_serial_rsci_ogwt & output_pxl_serial_rsci_irdy;
  assign output_pxl_serial_rsci_ogwt = output_pxl_serial_rsci_oswt & (~ output_pxl_serial_rsci_bcwt);
  assign output_pxl_serial_rsci_ivld_run_sct = output_pxl_serial_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_dp (
  clk, arst_n, atten_chan_out_rsci_oswt, atten_chan_out_rsci_wen_comp, atten_chan_out_rsci_biwt,
      atten_chan_out_rsci_bdwt, atten_chan_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input atten_chan_out_rsci_oswt;
  output atten_chan_out_rsci_wen_comp;
  input atten_chan_out_rsci_biwt;
  input atten_chan_out_rsci_bdwt;
  output atten_chan_out_rsci_bcwt;
  reg atten_chan_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign atten_chan_out_rsci_wen_comp = (~ atten_chan_out_rsci_oswt) | atten_chan_out_rsci_biwt
      | atten_chan_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      atten_chan_out_rsci_bcwt <= 1'b0;
    end
    else begin
      atten_chan_out_rsci_bcwt <= ~((~(atten_chan_out_rsci_bcwt | atten_chan_out_rsci_biwt))
          | atten_chan_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_ctrl
    (
  run_wen, atten_chan_out_rsci_oswt, atten_chan_out_rsci_irdy, atten_chan_out_rsci_biwt,
      atten_chan_out_rsci_bdwt, atten_chan_out_rsci_bcwt, atten_chan_out_rsci_ivld_run_sct
);
  input run_wen;
  input atten_chan_out_rsci_oswt;
  input atten_chan_out_rsci_irdy;
  output atten_chan_out_rsci_biwt;
  output atten_chan_out_rsci_bdwt;
  input atten_chan_out_rsci_bcwt;
  output atten_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire atten_chan_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign atten_chan_out_rsci_bdwt = atten_chan_out_rsci_oswt & run_wen;
  assign atten_chan_out_rsci_biwt = atten_chan_out_rsci_ogwt & atten_chan_out_rsci_irdy;
  assign atten_chan_out_rsci_ogwt = atten_chan_out_rsci_oswt & (~ atten_chan_out_rsci_bcwt);
  assign atten_chan_out_rsci_ivld_run_sct = atten_chan_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_dp (
  clk, arst_n, color_chan_out_rsci_oswt, color_chan_out_rsci_wen_comp, color_chan_out_rsci_biwt,
      color_chan_out_rsci_bdwt, color_chan_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input color_chan_out_rsci_oswt;
  output color_chan_out_rsci_wen_comp;
  input color_chan_out_rsci_biwt;
  input color_chan_out_rsci_bdwt;
  output color_chan_out_rsci_bcwt;
  reg color_chan_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign color_chan_out_rsci_wen_comp = (~ color_chan_out_rsci_oswt) | color_chan_out_rsci_biwt
      | color_chan_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_chan_out_rsci_bcwt <= 1'b0;
    end
    else begin
      color_chan_out_rsci_bcwt <= ~((~(color_chan_out_rsci_bcwt | color_chan_out_rsci_biwt))
          | color_chan_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_ctrl
    (
  run_wen, color_chan_out_rsci_oswt, color_chan_out_rsci_irdy, color_chan_out_rsci_biwt,
      color_chan_out_rsci_bdwt, color_chan_out_rsci_bcwt, color_chan_out_rsci_ivld_run_sct
);
  input run_wen;
  input color_chan_out_rsci_oswt;
  input color_chan_out_rsci_irdy;
  output color_chan_out_rsci_biwt;
  output color_chan_out_rsci_bdwt;
  input color_chan_out_rsci_bcwt;
  output color_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire color_chan_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign color_chan_out_rsci_bdwt = color_chan_out_rsci_oswt & run_wen;
  assign color_chan_out_rsci_biwt = color_chan_out_rsci_ogwt & color_chan_out_rsci_irdy;
  assign color_chan_out_rsci_ogwt = color_chan_out_rsci_oswt & (~ color_chan_out_rsci_bcwt);
  assign color_chan_out_rsci_ivld_run_sct = color_chan_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_out_rsci_params_out_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_out_rsci_params_out_wait_dp (
  clk, arst_n, params_out_rsci_oswt, params_out_rsci_wen_comp, params_out_rsci_biwt,
      params_out_rsci_bdwt, params_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input params_out_rsci_oswt;
  output params_out_rsci_wen_comp;
  input params_out_rsci_biwt;
  input params_out_rsci_bdwt;
  output params_out_rsci_bcwt;
  reg params_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign params_out_rsci_wen_comp = (~ params_out_rsci_oswt) | params_out_rsci_biwt
      | params_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_out_rsci_bcwt <= 1'b0;
    end
    else begin
      params_out_rsci_bcwt <= ~((~(params_out_rsci_bcwt | params_out_rsci_biwt))
          | params_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_out_rsci_params_out_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_out_rsci_params_out_wait_ctrl (
  run_wen, params_out_rsci_oswt, params_out_rsci_irdy, params_out_rsci_biwt, params_out_rsci_bdwt,
      params_out_rsci_bcwt, params_out_rsci_ivld_run_sct
);
  input run_wen;
  input params_out_rsci_oswt;
  input params_out_rsci_irdy;
  output params_out_rsci_biwt;
  output params_out_rsci_bdwt;
  input params_out_rsci_bcwt;
  output params_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire params_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_out_rsci_bdwt = params_out_rsci_oswt & run_wen;
  assign params_out_rsci_biwt = params_out_rsci_ogwt & params_out_rsci_irdy;
  assign params_out_rsci_ogwt = params_out_rsci_oswt & (~ params_out_rsci_bcwt);
  assign params_out_rsci_ivld_run_sct = params_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_dp (
  clk, arst_n, ray_out_rsci_oswt, ray_out_rsci_wen_comp, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt
);
  input clk;
  input arst_n;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input ray_out_rsci_biwt;
  input ray_out_rsci_bdwt;
  output ray_out_rsci_bcwt;
  reg ray_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_wen_comp = (~ ray_out_rsci_oswt) | ray_out_rsci_biwt | ray_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_out_rsci_bcwt <= ~((~(ray_out_rsci_bcwt | ray_out_rsci_biwt)) | ray_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_ctrl (
  run_wen, ray_out_rsci_oswt, ray_out_rsci_irdy, ray_out_rsci_biwt, ray_out_rsci_bdwt,
      ray_out_rsci_bcwt, ray_out_rsci_ivld_run_sct
);
  input run_wen;
  input ray_out_rsci_oswt;
  input ray_out_rsci_irdy;
  output ray_out_rsci_biwt;
  output ray_out_rsci_bdwt;
  input ray_out_rsci_bcwt;
  output ray_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire ray_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_out_rsci_bdwt = ray_out_rsci_oswt & run_wen;
  assign ray_out_rsci_biwt = ray_out_rsci_ogwt & ray_out_rsci_irdy;
  assign ray_out_rsci_ogwt = ray_out_rsci_oswt & (~ ray_out_rsci_bcwt);
  assign ray_out_rsci_ivld_run_sct = ray_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_dp (
  clk, arst_n, atten_chan_in_rsci_oswt, atten_chan_in_rsci_wen_comp, atten_chan_in_rsci_idat_mxwt,
      atten_chan_in_rsci_biwt, atten_chan_in_rsci_bdwt, atten_chan_in_rsci_bcwt,
      atten_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input atten_chan_in_rsci_oswt;
  output atten_chan_in_rsci_wen_comp;
  output [80:0] atten_chan_in_rsci_idat_mxwt;
  input atten_chan_in_rsci_biwt;
  input atten_chan_in_rsci_bdwt;
  output atten_chan_in_rsci_bcwt;
  reg atten_chan_in_rsci_bcwt;
  input [80:0] atten_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] atten_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign atten_chan_in_rsci_wen_comp = (~ atten_chan_in_rsci_oswt) | atten_chan_in_rsci_biwt
      | atten_chan_in_rsci_bcwt;
  assign atten_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(atten_chan_in_rsci_idat, atten_chan_in_rsci_idat_bfwt,
      atten_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      atten_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      atten_chan_in_rsci_bcwt <= ~((~(atten_chan_in_rsci_bcwt | atten_chan_in_rsci_biwt))
          | atten_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      atten_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ atten_chan_in_rsci_bcwt ) begin
      atten_chan_in_rsci_idat_bfwt <= atten_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_ctrl (
  run_wen, atten_chan_in_rsci_oswt, atten_chan_in_rsci_biwt, atten_chan_in_rsci_bdwt,
      atten_chan_in_rsci_bcwt, atten_chan_in_rsci_irdy_run_sct, atten_chan_in_rsci_ivld
);
  input run_wen;
  input atten_chan_in_rsci_oswt;
  output atten_chan_in_rsci_biwt;
  output atten_chan_in_rsci_bdwt;
  input atten_chan_in_rsci_bcwt;
  output atten_chan_in_rsci_irdy_run_sct;
  input atten_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire atten_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign atten_chan_in_rsci_bdwt = atten_chan_in_rsci_oswt & run_wen;
  assign atten_chan_in_rsci_biwt = atten_chan_in_rsci_ogwt & atten_chan_in_rsci_ivld;
  assign atten_chan_in_rsci_ogwt = atten_chan_in_rsci_oswt & (~ atten_chan_in_rsci_bcwt);
  assign atten_chan_in_rsci_irdy_run_sct = atten_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_dp (
  clk, arst_n, color_chan_in_rsci_oswt, color_chan_in_rsci_wen_comp, color_chan_in_rsci_idat_mxwt,
      color_chan_in_rsci_biwt, color_chan_in_rsci_bdwt, color_chan_in_rsci_bcwt,
      color_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input color_chan_in_rsci_oswt;
  output color_chan_in_rsci_wen_comp;
  output [80:0] color_chan_in_rsci_idat_mxwt;
  input color_chan_in_rsci_biwt;
  input color_chan_in_rsci_bdwt;
  output color_chan_in_rsci_bcwt;
  reg color_chan_in_rsci_bcwt;
  input [80:0] color_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [80:0] color_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign color_chan_in_rsci_wen_comp = (~ color_chan_in_rsci_oswt) | color_chan_in_rsci_biwt
      | color_chan_in_rsci_bcwt;
  assign color_chan_in_rsci_idat_mxwt = MUX_v_81_2_2(color_chan_in_rsci_idat, color_chan_in_rsci_idat_bfwt,
      color_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      color_chan_in_rsci_bcwt <= ~((~(color_chan_in_rsci_bcwt | color_chan_in_rsci_biwt))
          | color_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_chan_in_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ color_chan_in_rsci_bcwt ) begin
      color_chan_in_rsci_idat_bfwt <= color_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_ctrl (
  run_wen, color_chan_in_rsci_oswt, color_chan_in_rsci_biwt, color_chan_in_rsci_bdwt,
      color_chan_in_rsci_bcwt, color_chan_in_rsci_irdy_run_sct, color_chan_in_rsci_ivld
);
  input run_wen;
  input color_chan_in_rsci_oswt;
  output color_chan_in_rsci_biwt;
  output color_chan_in_rsci_bdwt;
  input color_chan_in_rsci_bcwt;
  output color_chan_in_rsci_irdy_run_sct;
  input color_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire color_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign color_chan_in_rsci_bdwt = color_chan_in_rsci_oswt & run_wen;
  assign color_chan_in_rsci_biwt = color_chan_in_rsci_ogwt & color_chan_in_rsci_ivld;
  assign color_chan_in_rsci_ogwt = color_chan_in_rsci_oswt & (~ color_chan_in_rsci_bcwt);
  assign color_chan_in_rsci_irdy_run_sct = color_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_in_rsci_params_in_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_in_rsci_params_in_wait_dp (
  clk, arst_n, params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt,
      params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt, params_in_rsci_idat
);
  input clk;
  input arst_n;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [92:0] params_in_rsci_idat_mxwt;
  input params_in_rsci_biwt;
  input params_in_rsci_bdwt;
  output params_in_rsci_bcwt;
  reg params_in_rsci_bcwt;
  input [92:0] params_in_rsci_idat;


  // Interconnect Declarations
  reg [92:0] params_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_wen_comp = (~ params_in_rsci_oswt) | params_in_rsci_biwt
      | params_in_rsci_bcwt;
  assign params_in_rsci_idat_mxwt = MUX_v_93_2_2(params_in_rsci_idat, params_in_rsci_idat_bfwt,
      params_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_bcwt <= 1'b0;
    end
    else begin
      params_in_rsci_bcwt <= ~((~(params_in_rsci_bcwt | params_in_rsci_biwt)) | params_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_rsci_idat_bfwt <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ params_in_rsci_bcwt ) begin
      params_in_rsci_idat_bfwt <= params_in_rsci_idat_mxwt;
    end
  end

  function automatic [92:0] MUX_v_93_2_2;
    input [92:0] input_0;
    input [92:0] input_1;
    input [0:0] sel;
    reg [92:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_93_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_in_rsci_params_in_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_in_rsci_params_in_wait_ctrl (
  run_wen, params_in_rsci_oswt, params_in_rsci_biwt, params_in_rsci_bdwt, params_in_rsci_bcwt,
      params_in_rsci_irdy_run_sct, params_in_rsci_ivld
);
  input run_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_biwt;
  output params_in_rsci_bdwt;
  input params_in_rsci_bcwt;
  output params_in_rsci_irdy_run_sct;
  input params_in_rsci_ivld;


  // Interconnect Declarations
  wire params_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign params_in_rsci_bdwt = params_in_rsci_oswt & run_wen;
  assign params_in_rsci_biwt = params_in_rsci_ogwt & params_in_rsci_ivld;
  assign params_in_rsci_ogwt = params_in_rsci_oswt & (~ params_in_rsci_bcwt);
  assign params_in_rsci_irdy_run_sct = params_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_dp
    (
  clk, arst_n, ray_scattered_chan_rsci_oswt, ray_scattered_chan_rsci_wen_comp, ray_scattered_chan_rsci_idat_mxwt,
      ray_scattered_chan_rsci_biwt, ray_scattered_chan_rsci_bdwt, ray_scattered_chan_rsci_bcwt,
      ray_scattered_chan_rsci_idat
);
  input clk;
  input arst_n;
  input ray_scattered_chan_rsci_oswt;
  output ray_scattered_chan_rsci_wen_comp;
  output [165:0] ray_scattered_chan_rsci_idat_mxwt;
  input ray_scattered_chan_rsci_biwt;
  input ray_scattered_chan_rsci_bdwt;
  output ray_scattered_chan_rsci_bcwt;
  reg ray_scattered_chan_rsci_bcwt;
  input [165:0] ray_scattered_chan_rsci_idat;


  // Interconnect Declarations
  reg [165:0] ray_scattered_chan_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_scattered_chan_rsci_wen_comp = (~ ray_scattered_chan_rsci_oswt) | ray_scattered_chan_rsci_biwt
      | ray_scattered_chan_rsci_bcwt;
  assign ray_scattered_chan_rsci_idat_mxwt = MUX_v_166_2_2(ray_scattered_chan_rsci_idat,
      ray_scattered_chan_rsci_idat_bfwt, ray_scattered_chan_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_scattered_chan_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_scattered_chan_rsci_bcwt <= ~((~(ray_scattered_chan_rsci_bcwt | ray_scattered_chan_rsci_biwt))
          | ray_scattered_chan_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_scattered_chan_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_scattered_chan_rsci_bcwt ) begin
      ray_scattered_chan_rsci_idat_bfwt <= ray_scattered_chan_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_ctrl
    (
  run_wen, ray_scattered_chan_rsci_oswt, ray_scattered_chan_rsci_biwt, ray_scattered_chan_rsci_bdwt,
      ray_scattered_chan_rsci_bcwt, ray_scattered_chan_rsci_irdy_run_sct, ray_scattered_chan_rsci_ivld
);
  input run_wen;
  input ray_scattered_chan_rsci_oswt;
  output ray_scattered_chan_rsci_biwt;
  output ray_scattered_chan_rsci_bdwt;
  input ray_scattered_chan_rsci_bcwt;
  output ray_scattered_chan_rsci_irdy_run_sct;
  input ray_scattered_chan_rsci_ivld;


  // Interconnect Declarations
  wire ray_scattered_chan_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_scattered_chan_rsci_bdwt = ray_scattered_chan_rsci_oswt & run_wen;
  assign ray_scattered_chan_rsci_biwt = ray_scattered_chan_rsci_ogwt & ray_scattered_chan_rsci_ivld;
  assign ray_scattered_chan_rsci_ogwt = ray_scattered_chan_rsci_oswt & (~ ray_scattered_chan_rsci_bcwt);
  assign ray_scattered_chan_rsci_irdy_run_sct = ray_scattered_chan_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_dp
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_dp (
  clk, arst_n, ray_chan_in_rsci_oswt, ray_chan_in_rsci_wen_comp, ray_chan_in_rsci_idat_mxwt,
      ray_chan_in_rsci_biwt, ray_chan_in_rsci_bdwt, ray_chan_in_rsci_bcwt, ray_chan_in_rsci_idat
);
  input clk;
  input arst_n;
  input ray_chan_in_rsci_oswt;
  output ray_chan_in_rsci_wen_comp;
  output [165:0] ray_chan_in_rsci_idat_mxwt;
  input ray_chan_in_rsci_biwt;
  input ray_chan_in_rsci_bdwt;
  output ray_chan_in_rsci_bcwt;
  reg ray_chan_in_rsci_bcwt;
  input [165:0] ray_chan_in_rsci_idat;


  // Interconnect Declarations
  reg [165:0] ray_chan_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_chan_in_rsci_wen_comp = (~ ray_chan_in_rsci_oswt) | ray_chan_in_rsci_biwt
      | ray_chan_in_rsci_bcwt;
  assign ray_chan_in_rsci_idat_mxwt = MUX_v_166_2_2(ray_chan_in_rsci_idat, ray_chan_in_rsci_idat_bfwt,
      ray_chan_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_chan_in_rsci_bcwt <= 1'b0;
    end
    else begin
      ray_chan_in_rsci_bcwt <= ~((~(ray_chan_in_rsci_bcwt | ray_chan_in_rsci_biwt))
          | ray_chan_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_chan_in_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ ray_chan_in_rsci_bcwt ) begin
      ray_chan_in_rsci_idat_bfwt <= ray_chan_in_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_ctrl
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_ctrl (
  run_wen, ray_chan_in_rsci_oswt, ray_chan_in_rsci_biwt, ray_chan_in_rsci_bdwt, ray_chan_in_rsci_bcwt,
      ray_chan_in_rsci_irdy_run_sct, ray_chan_in_rsci_ivld
);
  input run_wen;
  input ray_chan_in_rsci_oswt;
  output ray_chan_in_rsci_biwt;
  output ray_chan_in_rsci_bdwt;
  input ray_chan_in_rsci_bcwt;
  output ray_chan_in_rsci_irdy_run_sct;
  input ray_chan_in_rsci_ivld;


  // Interconnect Declarations
  wire ray_chan_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ray_chan_in_rsci_bdwt = ray_chan_in_rsci_oswt & run_wen;
  assign ray_chan_in_rsci_biwt = ray_chan_in_rsci_ogwt & ray_chan_in_rsci_ivld;
  assign ray_chan_in_rsci_ogwt = ray_chan_in_rsci_oswt & (~ ray_chan_in_rsci_bcwt);
  assign ray_chan_in_rsci_irdy_run_sct = ray_chan_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module RayCollector_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, for_C_2_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input for_C_2_tr0;


  // FSM State Type Declaration for RayCollector_run_run_fsm_1
  parameter
    run_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    main_C_1 = 3'd2,
    for_C_0 = 3'd3,
    for_C_1 = 3'd4,
    for_C_2 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : RayCollector_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 6'b000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 6'b000100;
        state_var_NS = for_C_0;
      end
      for_C_0 : begin
        fsm_output = 6'b001000;
        state_var_NS = for_C_1;
      end
      for_C_1 : begin
        fsm_output = 6'b010000;
        state_var_NS = for_C_2;
      end
      for_C_2 : begin
        fsm_output = 6'b100000;
        if ( for_C_2_tr0 ) begin
          state_var_NS = main_C_0;
        end
        else begin
          state_var_NS = for_C_0;
        end
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 6'b000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_staller
// ------------------------------------------------------------------


module RayCollector_run_staller (
  run_wen, rayIn_rsci_wen_comp, paramsIn_rsci_wen_comp, paramsOut_rsci_wen_comp,
      rayOut_rsci_wen_comp
);
  output run_wen;
  input rayIn_rsci_wen_comp;
  input paramsIn_rsci_wen_comp;
  input paramsOut_rsci_wen_comp;
  input rayOut_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = rayIn_rsci_wen_comp & paramsIn_rsci_wen_comp & paramsOut_rsci_wen_comp
      & rayOut_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayOut_rsci_rayOut_wait_dp
// ------------------------------------------------------------------


module RayCollector_run_rayOut_rsci_rayOut_wait_dp (
  clk, arst_n, rayOut_rsci_oswt, rayOut_rsci_wen_comp, rayOut_rsci_biwt, rayOut_rsci_bdwt,
      rayOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input rayOut_rsci_oswt;
  output rayOut_rsci_wen_comp;
  input rayOut_rsci_biwt;
  input rayOut_rsci_bdwt;
  output rayOut_rsci_bcwt;
  reg rayOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rayOut_rsci_wen_comp = (~ rayOut_rsci_oswt) | rayOut_rsci_biwt | rayOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayOut_rsci_bcwt <= 1'b0;
    end
    else begin
      rayOut_rsci_bcwt <= ~((~(rayOut_rsci_bcwt | rayOut_rsci_biwt)) | rayOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayOut_rsci_rayOut_wait_ctrl
// ------------------------------------------------------------------


module RayCollector_run_rayOut_rsci_rayOut_wait_ctrl (
  run_wen, rayOut_rsci_oswt, rayOut_rsci_irdy, rayOut_rsci_biwt, rayOut_rsci_bdwt,
      rayOut_rsci_bcwt, rayOut_rsci_ivld_run_sct
);
  input run_wen;
  input rayOut_rsci_oswt;
  input rayOut_rsci_irdy;
  output rayOut_rsci_biwt;
  output rayOut_rsci_bdwt;
  input rayOut_rsci_bcwt;
  output rayOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire rayOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rayOut_rsci_bdwt = rayOut_rsci_oswt & run_wen;
  assign rayOut_rsci_biwt = rayOut_rsci_ogwt & rayOut_rsci_irdy;
  assign rayOut_rsci_ogwt = rayOut_rsci_oswt & (~ rayOut_rsci_bcwt);
  assign rayOut_rsci_ivld_run_sct = rayOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsOut_rsci_paramsOut_wait_dp
// ------------------------------------------------------------------


module RayCollector_run_paramsOut_rsci_paramsOut_wait_dp (
  clk, arst_n, paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_biwt,
      paramsOut_rsci_bdwt, paramsOut_rsci_bcwt
);
  input clk;
  input arst_n;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input paramsOut_rsci_biwt;
  input paramsOut_rsci_bdwt;
  output paramsOut_rsci_bcwt;
  reg paramsOut_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_wen_comp = (~ paramsOut_rsci_oswt) | paramsOut_rsci_biwt
      | paramsOut_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsOut_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsOut_rsci_bcwt <= ~((~(paramsOut_rsci_bcwt | paramsOut_rsci_biwt)) | paramsOut_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsOut_rsci_paramsOut_wait_ctrl
// ------------------------------------------------------------------


module RayCollector_run_paramsOut_rsci_paramsOut_wait_ctrl (
  run_wen, paramsOut_rsci_oswt, paramsOut_rsci_irdy, paramsOut_rsci_biwt, paramsOut_rsci_bdwt,
      paramsOut_rsci_bcwt, paramsOut_rsci_ivld_run_sct
);
  input run_wen;
  input paramsOut_rsci_oswt;
  input paramsOut_rsci_irdy;
  output paramsOut_rsci_biwt;
  output paramsOut_rsci_bdwt;
  input paramsOut_rsci_bcwt;
  output paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire paramsOut_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsOut_rsci_bdwt = paramsOut_rsci_oswt & run_wen;
  assign paramsOut_rsci_biwt = paramsOut_rsci_ogwt & paramsOut_rsci_irdy;
  assign paramsOut_rsci_ogwt = paramsOut_rsci_oswt & (~ paramsOut_rsci_bcwt);
  assign paramsOut_rsci_ivld_run_sct = paramsOut_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsIn_rsci_paramsIn_wait_dp
// ------------------------------------------------------------------


module RayCollector_run_paramsIn_rsci_paramsIn_wait_dp (
  clk, arst_n, paramsIn_rsci_oswt, paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt,
      paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt, paramsIn_rsci_idat
);
  input clk;
  input arst_n;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [92:0] paramsIn_rsci_idat_mxwt;
  input paramsIn_rsci_biwt;
  input paramsIn_rsci_bdwt;
  output paramsIn_rsci_bcwt;
  reg paramsIn_rsci_bcwt;
  input [92:0] paramsIn_rsci_idat;


  // Interconnect Declarations
  reg [92:0] paramsIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_wen_comp = (~ paramsIn_rsci_oswt) | paramsIn_rsci_biwt | paramsIn_rsci_bcwt;
  assign paramsIn_rsci_idat_mxwt = MUX_v_93_2_2(paramsIn_rsci_idat, paramsIn_rsci_idat_bfwt,
      paramsIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_bcwt <= 1'b0;
    end
    else begin
      paramsIn_rsci_bcwt <= ~((~(paramsIn_rsci_bcwt | paramsIn_rsci_biwt)) | paramsIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_rsci_idat_bfwt <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ paramsIn_rsci_bcwt ) begin
      paramsIn_rsci_idat_bfwt <= paramsIn_rsci_idat_mxwt;
    end
  end

  function automatic [92:0] MUX_v_93_2_2;
    input [92:0] input_0;
    input [92:0] input_1;
    input [0:0] sel;
    reg [92:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_93_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsIn_rsci_paramsIn_wait_ctrl
// ------------------------------------------------------------------


module RayCollector_run_paramsIn_rsci_paramsIn_wait_ctrl (
  run_wen, paramsIn_rsci_oswt, paramsIn_rsci_biwt, paramsIn_rsci_bdwt, paramsIn_rsci_bcwt,
      paramsIn_rsci_irdy_run_sct, paramsIn_rsci_ivld
);
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_biwt;
  output paramsIn_rsci_bdwt;
  input paramsIn_rsci_bcwt;
  output paramsIn_rsci_irdy_run_sct;
  input paramsIn_rsci_ivld;


  // Interconnect Declarations
  wire paramsIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign paramsIn_rsci_bdwt = paramsIn_rsci_oswt & run_wen;
  assign paramsIn_rsci_biwt = paramsIn_rsci_ogwt & paramsIn_rsci_ivld;
  assign paramsIn_rsci_ogwt = paramsIn_rsci_oswt & (~ paramsIn_rsci_bcwt);
  assign paramsIn_rsci_irdy_run_sct = paramsIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayIn_rsci_rayIn_wait_dp
// ------------------------------------------------------------------


module RayCollector_run_rayIn_rsci_rayIn_wait_dp (
  clk, arst_n, rayIn_rsci_oswt, rayIn_rsci_wen_comp, rayIn_rsci_idat_mxwt, rayIn_rsci_biwt,
      rayIn_rsci_bdwt, rayIn_rsci_bcwt, rayIn_rsci_idat
);
  input clk;
  input arst_n;
  input rayIn_rsci_oswt;
  output rayIn_rsci_wen_comp;
  output [165:0] rayIn_rsci_idat_mxwt;
  input rayIn_rsci_biwt;
  input rayIn_rsci_bdwt;
  output rayIn_rsci_bcwt;
  reg rayIn_rsci_bcwt;
  input [165:0] rayIn_rsci_idat;


  // Interconnect Declarations
  reg [165:0] rayIn_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rayIn_rsci_wen_comp = (~ rayIn_rsci_oswt) | rayIn_rsci_biwt | rayIn_rsci_bcwt;
  assign rayIn_rsci_idat_mxwt = MUX_v_166_2_2(rayIn_rsci_idat, rayIn_rsci_idat_bfwt,
      rayIn_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayIn_rsci_bcwt <= 1'b0;
    end
    else begin
      rayIn_rsci_bcwt <= ~((~(rayIn_rsci_bcwt | rayIn_rsci_biwt)) | rayIn_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayIn_rsci_idat_bfwt <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ rayIn_rsci_bcwt ) begin
      rayIn_rsci_idat_bfwt <= rayIn_rsci_idat_mxwt;
    end
  end

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayIn_rsci_rayIn_wait_ctrl
// ------------------------------------------------------------------


module RayCollector_run_rayIn_rsci_rayIn_wait_ctrl (
  run_wen, rayIn_rsci_oswt, rayIn_rsci_biwt, rayIn_rsci_bdwt, rayIn_rsci_bcwt, rayIn_rsci_irdy_run_sct,
      rayIn_rsci_ivld
);
  input run_wen;
  input rayIn_rsci_oswt;
  output rayIn_rsci_biwt;
  output rayIn_rsci_bdwt;
  input rayIn_rsci_bcwt;
  output rayIn_rsci_irdy_run_sct;
  input rayIn_rsci_ivld;


  // Interconnect Declarations
  wire rayIn_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign rayIn_rsci_bdwt = rayIn_rsci_oswt & run_wen;
  assign rayIn_rsci_biwt = rayIn_rsci_ogwt & rayIn_rsci_ivld;
  assign rayIn_rsci_ogwt = rayIn_rsci_oswt & (~ rayIn_rsci_bcwt);
  assign rayIn_rsci_irdy_run_sct = rayIn_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_staller
// ------------------------------------------------------------------


module PixelAccumulator_run_staller (
  run_wen, accumulator_parms_rsci_wen_comp, pxl_sample_rsci_wen_comp, output_pxl_serial_rsci_wen_comp
);
  output run_wen;
  input accumulator_parms_rsci_wen_comp;
  input pxl_sample_rsci_wen_comp;
  input output_pxl_serial_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = accumulator_parms_rsci_wen_comp & pxl_sample_rsci_wen_comp & output_pxl_serial_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp
// ------------------------------------------------------------------


module PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp (
  clk, arst_n, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_wen_comp, output_pxl_serial_rsci_biwt,
      output_pxl_serial_rsci_bdwt, output_pxl_serial_rsci_bcwt
);
  input clk;
  input arst_n;
  input output_pxl_serial_rsci_oswt;
  output output_pxl_serial_rsci_wen_comp;
  input output_pxl_serial_rsci_biwt;
  input output_pxl_serial_rsci_bdwt;
  output output_pxl_serial_rsci_bcwt;
  reg output_pxl_serial_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign output_pxl_serial_rsci_wen_comp = (~ output_pxl_serial_rsci_oswt) | output_pxl_serial_rsci_biwt
      | output_pxl_serial_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_pxl_serial_rsci_bcwt <= 1'b0;
    end
    else begin
      output_pxl_serial_rsci_bcwt <= ~((~(output_pxl_serial_rsci_bcwt | output_pxl_serial_rsci_biwt))
          | output_pxl_serial_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl
// ------------------------------------------------------------------


module PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl (
  run_wen, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_irdy, output_pxl_serial_rsci_biwt,
      output_pxl_serial_rsci_bdwt, output_pxl_serial_rsci_bcwt, output_pxl_serial_rsci_ivld_run_sct
);
  input run_wen;
  input output_pxl_serial_rsci_oswt;
  input output_pxl_serial_rsci_irdy;
  output output_pxl_serial_rsci_biwt;
  output output_pxl_serial_rsci_bdwt;
  input output_pxl_serial_rsci_bcwt;
  output output_pxl_serial_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire output_pxl_serial_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign output_pxl_serial_rsci_bdwt = output_pxl_serial_rsci_oswt & run_wen;
  assign output_pxl_serial_rsci_biwt = output_pxl_serial_rsci_ogwt & output_pxl_serial_rsci_irdy;
  assign output_pxl_serial_rsci_ogwt = output_pxl_serial_rsci_oswt & (~ output_pxl_serial_rsci_bcwt);
  assign output_pxl_serial_rsci_ivld_run_sct = output_pxl_serial_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_dp
// ------------------------------------------------------------------


module PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_dp (
  clk, arst_n, pxl_sample_rsci_oswt, pxl_sample_rsci_wen_comp, pxl_sample_rsci_idat_mxwt,
      pxl_sample_rsci_biwt, pxl_sample_rsci_bdwt, pxl_sample_rsci_bcwt, pxl_sample_rsci_idat
);
  input clk;
  input arst_n;
  input pxl_sample_rsci_oswt;
  output pxl_sample_rsci_wen_comp;
  output [80:0] pxl_sample_rsci_idat_mxwt;
  input pxl_sample_rsci_biwt;
  input pxl_sample_rsci_bdwt;
  output pxl_sample_rsci_bcwt;
  reg pxl_sample_rsci_bcwt;
  input [80:0] pxl_sample_rsci_idat;


  // Interconnect Declarations
  reg [80:0] pxl_sample_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign pxl_sample_rsci_wen_comp = (~ pxl_sample_rsci_oswt) | pxl_sample_rsci_biwt
      | pxl_sample_rsci_bcwt;
  assign pxl_sample_rsci_idat_mxwt = MUX_v_81_2_2(pxl_sample_rsci_idat, pxl_sample_rsci_idat_bfwt,
      pxl_sample_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pxl_sample_rsci_bcwt <= 1'b0;
    end
    else begin
      pxl_sample_rsci_bcwt <= ~((~(pxl_sample_rsci_bcwt | pxl_sample_rsci_biwt))
          | pxl_sample_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pxl_sample_rsci_idat_bfwt <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ pxl_sample_rsci_bcwt ) begin
      pxl_sample_rsci_idat_bfwt <= pxl_sample_rsci_idat_mxwt;
    end
  end

  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_ctrl
// ------------------------------------------------------------------


module PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_ctrl (
  run_wen, pxl_sample_rsci_oswt, pxl_sample_rsci_biwt, pxl_sample_rsci_bdwt, pxl_sample_rsci_bcwt,
      pxl_sample_rsci_irdy_run_sct, pxl_sample_rsci_ivld
);
  input run_wen;
  input pxl_sample_rsci_oswt;
  output pxl_sample_rsci_biwt;
  output pxl_sample_rsci_bdwt;
  input pxl_sample_rsci_bcwt;
  output pxl_sample_rsci_irdy_run_sct;
  input pxl_sample_rsci_ivld;


  // Interconnect Declarations
  wire pxl_sample_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign pxl_sample_rsci_bdwt = pxl_sample_rsci_oswt & run_wen;
  assign pxl_sample_rsci_biwt = pxl_sample_rsci_ogwt & pxl_sample_rsci_ivld;
  assign pxl_sample_rsci_ogwt = pxl_sample_rsci_oswt & (~ pxl_sample_rsci_bcwt);
  assign pxl_sample_rsci_irdy_run_sct = pxl_sample_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_dp
// ------------------------------------------------------------------


module PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_dp (
  clk, arst_n, accumulator_parms_rsci_oswt, accumulator_parms_rsci_wen_comp, accumulator_parms_rsci_idat_mxwt,
      accumulator_parms_rsci_biwt, accumulator_parms_rsci_bdwt, accumulator_parms_rsci_bcwt,
      accumulator_parms_rsci_idat
);
  input clk;
  input arst_n;
  input accumulator_parms_rsci_oswt;
  output accumulator_parms_rsci_wen_comp;
  output [34:0] accumulator_parms_rsci_idat_mxwt;
  input accumulator_parms_rsci_biwt;
  input accumulator_parms_rsci_bdwt;
  output accumulator_parms_rsci_bcwt;
  reg accumulator_parms_rsci_bcwt;
  input [419:0] accumulator_parms_rsci_idat;


  // Interconnect Declarations
  reg [32:0] reg_accumulator_parms_rsci_idat_bfwt_ftd;
  reg [1:0] reg_accumulator_parms_rsci_idat_bfwt_ftd_93;
  wire [32:0] accumulator_parms_rsci_idat_mxwt_opt_137_105;
  wire [1:0] accumulator_parms_rsci_idat_mxwt_opt_12_11;


  // Interconnect Declarations for Component Instantiations 
  assign accumulator_parms_rsci_wen_comp = (~ accumulator_parms_rsci_oswt) | accumulator_parms_rsci_biwt
      | accumulator_parms_rsci_bcwt;
  assign accumulator_parms_rsci_idat_mxwt_opt_137_105 = MUX_v_33_2_2((accumulator_parms_rsci_idat[137:105]),
      reg_accumulator_parms_rsci_idat_bfwt_ftd, accumulator_parms_rsci_bcwt);
  assign accumulator_parms_rsci_idat_mxwt_opt_12_11 = MUX_v_2_2_2((accumulator_parms_rsci_idat[12:11]),
      reg_accumulator_parms_rsci_idat_bfwt_ftd_93, accumulator_parms_rsci_bcwt);
  assign accumulator_parms_rsci_idat_mxwt = {accumulator_parms_rsci_idat_mxwt_opt_137_105
      , accumulator_parms_rsci_idat_mxwt_opt_12_11};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulator_parms_rsci_bcwt <= 1'b0;
    end
    else begin
      accumulator_parms_rsci_bcwt <= ~((~(accumulator_parms_rsci_bcwt | accumulator_parms_rsci_biwt))
          | accumulator_parms_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_accumulator_parms_rsci_idat_bfwt_ftd <= 33'b000000000000000000000000000000000;
    end
    else if ( ~ accumulator_parms_rsci_bcwt ) begin
      reg_accumulator_parms_rsci_idat_bfwt_ftd <= accumulator_parms_rsci_idat_mxwt_opt_137_105;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_accumulator_parms_rsci_idat_bfwt_ftd_93 <= 2'b00;
    end
    else if ( ~ accumulator_parms_rsci_bcwt ) begin
      reg_accumulator_parms_rsci_idat_bfwt_ftd_93 <= accumulator_parms_rsci_idat_mxwt_opt_12_11;
    end
  end

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [32:0] MUX_v_33_2_2;
    input [32:0] input_0;
    input [32:0] input_1;
    input [0:0] sel;
    reg [32:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_33_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_ctrl
// ------------------------------------------------------------------


module PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_ctrl (
  run_wen, accumulator_parms_rsci_oswt, accumulator_parms_rsci_biwt, accumulator_parms_rsci_bdwt,
      accumulator_parms_rsci_bcwt, accumulator_parms_rsci_irdy_run_sct, accumulator_parms_rsci_ivld
);
  input run_wen;
  input accumulator_parms_rsci_oswt;
  output accumulator_parms_rsci_biwt;
  output accumulator_parms_rsci_bdwt;
  input accumulator_parms_rsci_bcwt;
  output accumulator_parms_rsci_irdy_run_sct;
  input accumulator_parms_rsci_ivld;


  // Interconnect Declarations
  wire accumulator_parms_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign accumulator_parms_rsci_bdwt = accumulator_parms_rsci_oswt & run_wen;
  assign accumulator_parms_rsci_biwt = accumulator_parms_rsci_ogwt & accumulator_parms_rsci_ivld;
  assign accumulator_parms_rsci_ogwt = accumulator_parms_rsci_oswt & (~ accumulator_parms_rsci_bcwt);
  assign accumulator_parms_rsci_irdy_run_sct = accumulator_parms_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_quad_serial_out_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_quad_serial_out_rsci (
  clk, arst_n, quad_serial_out_rsc_dat, quad_serial_out_rsc_vld, quad_serial_out_rsc_rdy,
      run_wen, quad_serial_out_rsci_oswt, quad_serial_out_rsci_wen_comp, quad_serial_out_rsci_idat
);
  input clk;
  input arst_n;
  output [376:0] quad_serial_out_rsc_dat;
  output quad_serial_out_rsc_vld;
  input quad_serial_out_rsc_rdy;
  input run_wen;
  input quad_serial_out_rsci_oswt;
  output quad_serial_out_rsci_wen_comp;
  input [376:0] quad_serial_out_rsci_idat;


  // Interconnect Declarations
  wire quad_serial_out_rsci_irdy;
  wire quad_serial_out_rsci_biwt;
  wire quad_serial_out_rsci_bdwt;
  wire quad_serial_out_rsci_bcwt;
  wire quad_serial_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd5),
  .width(32'sd377)) quad_serial_out_rsci (
      .irdy(quad_serial_out_rsci_irdy),
      .ivld(quad_serial_out_rsci_ivld_run_sct),
      .idat(quad_serial_out_rsci_idat),
      .rdy(quad_serial_out_rsc_rdy),
      .vld(quad_serial_out_rsc_vld),
      .dat(quad_serial_out_rsc_dat)
    );
  ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_ctrl ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quad_serial_out_rsci_oswt(quad_serial_out_rsci_oswt),
      .quad_serial_out_rsci_irdy(quad_serial_out_rsci_irdy),
      .quad_serial_out_rsci_biwt(quad_serial_out_rsci_biwt),
      .quad_serial_out_rsci_bdwt(quad_serial_out_rsci_bdwt),
      .quad_serial_out_rsci_bcwt(quad_serial_out_rsci_bcwt),
      .quad_serial_out_rsci_ivld_run_sct(quad_serial_out_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_dp ParamsDeserializer_run_quad_serial_out_rsci_quad_serial_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_serial_out_rsci_oswt(quad_serial_out_rsci_oswt),
      .quad_serial_out_rsci_wen_comp(quad_serial_out_rsci_wen_comp),
      .quad_serial_out_rsci_biwt(quad_serial_out_rsci_biwt),
      .quad_serial_out_rsci_bdwt(quad_serial_out_rsci_bdwt),
      .quad_serial_out_rsci_bcwt(quad_serial_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_accum_params_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_accum_params_rsci (
  clk, arst_n, accum_params_rsc_dat, accum_params_rsc_vld, accum_params_rsc_rdy,
      run_wen, accum_params_rsci_oswt, accum_params_rsci_wen_comp, accum_params_rsci_idat
);
  input clk;
  input arst_n;
  output [419:0] accum_params_rsc_dat;
  output accum_params_rsc_vld;
  input accum_params_rsc_rdy;
  input run_wen;
  input accum_params_rsci_oswt;
  output accum_params_rsci_wen_comp;
  input [419:0] accum_params_rsci_idat;


  // Interconnect Declarations
  wire accum_params_rsci_irdy;
  wire accum_params_rsci_biwt;
  wire accum_params_rsci_bdwt;
  wire accum_params_rsci_bcwt;
  wire accum_params_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd4),
  .width(32'sd420)) accum_params_rsci (
      .irdy(accum_params_rsci_irdy),
      .ivld(accum_params_rsci_ivld_run_sct),
      .idat(accum_params_rsci_idat),
      .rdy(accum_params_rsc_rdy),
      .vld(accum_params_rsc_vld),
      .dat(accum_params_rsc_dat)
    );
  ParamsDeserializer_run_accum_params_rsci_accum_params_wait_ctrl ParamsDeserializer_run_accum_params_rsci_accum_params_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .accum_params_rsci_oswt(accum_params_rsci_oswt),
      .accum_params_rsci_irdy(accum_params_rsci_irdy),
      .accum_params_rsci_biwt(accum_params_rsci_biwt),
      .accum_params_rsci_bdwt(accum_params_rsci_bdwt),
      .accum_params_rsci_bcwt(accum_params_rsci_bcwt),
      .accum_params_rsci_ivld_run_sct(accum_params_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_accum_params_rsci_accum_params_wait_dp ParamsDeserializer_run_accum_params_rsci_accum_params_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accum_params_rsci_oswt(accum_params_rsci_oswt),
      .accum_params_rsci_wen_comp(accum_params_rsci_wen_comp),
      .accum_params_rsci_biwt(accum_params_rsci_biwt),
      .accum_params_rsci_bdwt(accum_params_rsci_bdwt),
      .accum_params_rsci_bcwt(accum_params_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_render_params_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_render_params_rsci (
  clk, arst_n, render_params_rsc_dat, render_params_rsc_vld, render_params_rsc_rdy,
      run_wen, render_params_rsci_oswt, render_params_rsci_wen_comp, render_params_rsci_idat
);
  input clk;
  input arst_n;
  output [419:0] render_params_rsc_dat;
  output render_params_rsc_vld;
  input render_params_rsc_rdy;
  input run_wen;
  input render_params_rsci_oswt;
  output render_params_rsci_wen_comp;
  input [419:0] render_params_rsci_idat;


  // Interconnect Declarations
  wire render_params_rsci_irdy;
  wire render_params_rsci_biwt;
  wire render_params_rsci_bdwt;
  wire render_params_rsci_bcwt;
  wire render_params_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd420)) render_params_rsci (
      .irdy(render_params_rsci_irdy),
      .ivld(render_params_rsci_ivld_run_sct),
      .idat(render_params_rsci_idat),
      .rdy(render_params_rsc_rdy),
      .vld(render_params_rsc_vld),
      .dat(render_params_rsc_dat)
    );
  ParamsDeserializer_run_render_params_rsci_render_params_wait_ctrl ParamsDeserializer_run_render_params_rsci_render_params_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .render_params_rsci_oswt(render_params_rsci_oswt),
      .render_params_rsci_irdy(render_params_rsci_irdy),
      .render_params_rsci_biwt(render_params_rsci_biwt),
      .render_params_rsci_bdwt(render_params_rsci_bdwt),
      .render_params_rsci_bcwt(render_params_rsci_bcwt),
      .render_params_rsci_ivld_run_sct(render_params_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_render_params_rsci_render_params_wait_dp ParamsDeserializer_run_render_params_rsci_render_params_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsci_oswt(render_params_rsci_oswt),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .render_params_rsci_biwt(render_params_rsci_biwt),
      .render_params_rsci_bdwt(render_params_rsci_bdwt),
      .render_params_rsci_bcwt(render_params_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_qbuffer_params_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_qbuffer_params_rsci (
  clk, arst_n, qbuffer_params_rsc_dat, qbuffer_params_rsc_vld, qbuffer_params_rsc_rdy,
      run_wen, qbuffer_params_rsci_oswt, qbuffer_params_rsci_wen_comp, qbuffer_params_rsci_idat
);
  input clk;
  input arst_n;
  output [56:0] qbuffer_params_rsc_dat;
  output qbuffer_params_rsc_vld;
  input qbuffer_params_rsc_rdy;
  input run_wen;
  input qbuffer_params_rsci_oswt;
  output qbuffer_params_rsci_wen_comp;
  input [56:0] qbuffer_params_rsci_idat;


  // Interconnect Declarations
  wire qbuffer_params_rsci_irdy;
  wire qbuffer_params_rsci_biwt;
  wire qbuffer_params_rsci_bdwt;
  wire qbuffer_params_rsci_bcwt;
  wire qbuffer_params_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd2),
  .width(32'sd57)) qbuffer_params_rsci (
      .irdy(qbuffer_params_rsci_irdy),
      .ivld(qbuffer_params_rsci_ivld_run_sct),
      .idat(qbuffer_params_rsci_idat),
      .rdy(qbuffer_params_rsc_rdy),
      .vld(qbuffer_params_rsc_vld),
      .dat(qbuffer_params_rsc_dat)
    );
  ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_ctrl ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .qbuffer_params_rsci_oswt(qbuffer_params_rsci_oswt),
      .qbuffer_params_rsci_irdy(qbuffer_params_rsci_irdy),
      .qbuffer_params_rsci_biwt(qbuffer_params_rsci_biwt),
      .qbuffer_params_rsci_bdwt(qbuffer_params_rsci_bdwt),
      .qbuffer_params_rsci_bcwt(qbuffer_params_rsci_bcwt),
      .qbuffer_params_rsci_ivld_run_sct(qbuffer_params_rsci_ivld_run_sct)
    );
  ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_dp ParamsDeserializer_run_qbuffer_params_rsci_qbuffer_params_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .qbuffer_params_rsci_oswt(qbuffer_params_rsci_oswt),
      .qbuffer_params_rsci_wen_comp(qbuffer_params_rsci_wen_comp),
      .qbuffer_params_rsci_biwt(qbuffer_params_rsci_biwt),
      .qbuffer_params_rsci_bdwt(qbuffer_params_rsci_bdwt),
      .qbuffer_params_rsci_bcwt(qbuffer_params_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run_inputChannel_rsci
// ------------------------------------------------------------------


module ParamsDeserializer_run_inputChannel_rsci (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      run_wen, inputChannel_rsci_oswt, inputChannel_rsci_wen_comp, inputChannel_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [11:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  input run_wen;
  input inputChannel_rsci_oswt;
  output inputChannel_rsci_wen_comp;
  output [11:0] inputChannel_rsci_idat_mxwt;


  // Interconnect Declarations
  wire inputChannel_rsci_biwt;
  wire inputChannel_rsci_bdwt;
  wire inputChannel_rsci_bcwt;
  wire inputChannel_rsci_irdy_run_sct;
  wire inputChannel_rsci_ivld;
  wire [11:0] inputChannel_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd12)) inputChannel_rsci (
      .rdy(inputChannel_rsc_rdy),
      .vld(inputChannel_rsc_vld),
      .dat(inputChannel_rsc_dat),
      .irdy(inputChannel_rsci_irdy_run_sct),
      .ivld(inputChannel_rsci_ivld),
      .idat(inputChannel_rsci_idat)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_irdy_run_sct(inputChannel_rsci_irdy_run_sct),
      .inputChannel_rsci_ivld(inputChannel_rsci_ivld)
    );
  ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp ParamsDeserializer_run_inputChannel_rsci_inputChannel_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsci_oswt(inputChannel_rsci_oswt),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt),
      .inputChannel_rsci_biwt(inputChannel_rsci_biwt),
      .inputChannel_rsci_bdwt(inputChannel_rsci_bdwt),
      .inputChannel_rsci_bcwt(inputChannel_rsci_bcwt),
      .inputChannel_rsci_idat(inputChannel_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_out_rsci
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_out_rsci (
  clk, arst_n, quads_out_rsc_dat, quads_out_rsc_vld, quads_out_rsc_rdy, run_wen,
      quads_out_rsci_oswt, quads_out_rsci_wen_comp, quads_out_rsci_idat
);
  input clk;
  input arst_n;
  output [376:0] quads_out_rsc_dat;
  output quads_out_rsc_vld;
  input quads_out_rsc_rdy;
  input run_wen;
  input quads_out_rsci_oswt;
  output quads_out_rsci_wen_comp;
  input [376:0] quads_out_rsci_idat;


  // Interconnect Declarations
  wire quads_out_rsci_irdy;
  wire quads_out_rsci_biwt;
  wire quads_out_rsci_bdwt;
  wire quads_out_rsci_bcwt;
  wire quads_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd377)) quads_out_rsci (
      .irdy(quads_out_rsci_irdy),
      .ivld(quads_out_rsci_ivld_run_sct),
      .idat(quads_out_rsci_idat),
      .rdy(quads_out_rsc_rdy),
      .vld(quads_out_rsc_vld),
      .dat(quads_out_rsc_dat)
    );
  QuadBuffer_64_run_quads_out_rsci_quads_out_wait_ctrl QuadBuffer_64_run_quads_out_rsci_quads_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quads_out_rsci_oswt(quads_out_rsci_oswt),
      .quads_out_rsci_irdy(quads_out_rsci_irdy),
      .quads_out_rsci_biwt(quads_out_rsci_biwt),
      .quads_out_rsci_bdwt(quads_out_rsci_bdwt),
      .quads_out_rsci_bcwt(quads_out_rsci_bcwt),
      .quads_out_rsci_ivld_run_sct(quads_out_rsci_ivld_run_sct)
    );
  QuadBuffer_64_run_quads_out_rsci_quads_out_wait_dp QuadBuffer_64_run_quads_out_rsci_quads_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quads_out_rsci_oswt(quads_out_rsci_oswt),
      .quads_out_rsci_wen_comp(quads_out_rsci_wen_comp),
      .quads_out_rsci_biwt(quads_out_rsci_biwt),
      .quads_out_rsci_bdwt(quads_out_rsci_bdwt),
      .quads_out_rsci_bcwt(quads_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_paramsIn_rsci
// ------------------------------------------------------------------


module QuadBuffer_64_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [56:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [45:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [56:0] paramsIn_rsci_idat;
  wire [45:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd7),
  .width(32'sd57)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_ctrl QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_dp QuadBuffer_64_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run_quads_in_rsci
// ------------------------------------------------------------------


module QuadBuffer_64_run_quads_in_rsci (
  clk, arst_n, quads_in_rsc_dat, quads_in_rsc_vld, quads_in_rsc_rdy, run_wen, quads_in_rsci_oswt,
      quads_in_rsci_wen_comp, quads_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [376:0] quads_in_rsc_dat;
  input quads_in_rsc_vld;
  output quads_in_rsc_rdy;
  input run_wen;
  input quads_in_rsci_oswt;
  output quads_in_rsci_wen_comp;
  output [376:0] quads_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quads_in_rsci_biwt;
  wire quads_in_rsci_bdwt;
  wire quads_in_rsci_bcwt;
  wire quads_in_rsci_irdy_run_sct;
  wire quads_in_rsci_ivld;
  wire [376:0] quads_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd377)) quads_in_rsci (
      .rdy(quads_in_rsc_rdy),
      .vld(quads_in_rsc_vld),
      .dat(quads_in_rsc_dat),
      .irdy(quads_in_rsci_irdy_run_sct),
      .ivld(quads_in_rsci_ivld),
      .idat(quads_in_rsci_idat)
    );
  QuadBuffer_64_run_quads_in_rsci_quads_in_wait_ctrl QuadBuffer_64_run_quads_in_rsci_quads_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quads_in_rsci_oswt(quads_in_rsci_oswt),
      .quads_in_rsci_biwt(quads_in_rsci_biwt),
      .quads_in_rsci_bdwt(quads_in_rsci_bdwt),
      .quads_in_rsci_bcwt(quads_in_rsci_bcwt),
      .quads_in_rsci_irdy_run_sct(quads_in_rsci_irdy_run_sct),
      .quads_in_rsci_ivld(quads_in_rsci_ivld)
    );
  QuadBuffer_64_run_quads_in_rsci_quads_in_wait_dp QuadBuffer_64_run_quads_in_rsci_quads_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsci_oswt(quads_in_rsci_oswt),
      .quads_in_rsci_wen_comp(quads_in_rsci_wen_comp),
      .quads_in_rsci_idat_mxwt(quads_in_rsci_idat_mxwt),
      .quads_in_rsci_biwt(quads_in_rsci_biwt),
      .quads_in_rsci_bdwt(quads_in_rsci_bdwt),
      .quads_in_rsci_bcwt(quads_in_rsci_bcwt),
      .quads_in_rsci_idat(quads_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_loopIndicesOut_rsci
// ------------------------------------------------------------------


module RenderLooper_run_loopIndicesOut_rsci (
  clk, arst_n, loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld, loopIndicesOut_rsc_rdy,
      run_wen, loopIndicesOut_rsci_oswt, loopIndicesOut_rsci_wen_comp, loopIndicesOut_rsci_idat
);
  input clk;
  input arst_n;
  output [22:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;
  input run_wen;
  input loopIndicesOut_rsci_oswt;
  output loopIndicesOut_rsci_wen_comp;
  input [22:0] loopIndicesOut_rsci_idat;


  // Interconnect Declarations
  wire loopIndicesOut_rsci_irdy;
  wire loopIndicesOut_rsci_biwt;
  wire loopIndicesOut_rsci_bdwt;
  wire loopIndicesOut_rsci_bcwt;
  wire loopIndicesOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd23),
  .width(32'sd23)) loopIndicesOut_rsci (
      .irdy(loopIndicesOut_rsci_irdy),
      .ivld(loopIndicesOut_rsci_ivld_run_sct),
      .idat(loopIndicesOut_rsci_idat),
      .rdy(loopIndicesOut_rsc_rdy),
      .vld(loopIndicesOut_rsc_vld),
      .dat(loopIndicesOut_rsc_dat)
    );
  RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_irdy(loopIndicesOut_rsci_irdy),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt),
      .loopIndicesOut_rsci_ivld_run_sct(loopIndicesOut_rsci_ivld_run_sct)
    );
  RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp RenderLooper_run_loopIndicesOut_rsci_loopIndicesOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsci_oswt(loopIndicesOut_rsci_oswt),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_biwt(loopIndicesOut_rsci_biwt),
      .loopIndicesOut_rsci_bdwt(loopIndicesOut_rsci_bdwt),
      .loopIndicesOut_rsci_bcwt(loopIndicesOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_out_rsci
// ------------------------------------------------------------------


module RenderLooper_run_render_params_out_rsci (
  clk, arst_n, render_params_out_rsc_dat, render_params_out_rsc_vld, render_params_out_rsc_rdy,
      run_wen, render_params_out_rsci_oswt, render_params_out_rsci_wen_comp, render_params_out_rsci_idat
);
  input clk;
  input arst_n;
  output [419:0] render_params_out_rsc_dat;
  output render_params_out_rsc_vld;
  input render_params_out_rsc_rdy;
  input run_wen;
  input render_params_out_rsci_oswt;
  output render_params_out_rsci_wen_comp;
  input [419:0] render_params_out_rsci_idat;


  // Interconnect Declarations
  wire render_params_out_rsci_irdy;
  wire render_params_out_rsci_biwt;
  wire render_params_out_rsci_bdwt;
  wire render_params_out_rsci_bcwt;
  wire render_params_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd22),
  .width(32'sd420)) render_params_out_rsci (
      .irdy(render_params_out_rsci_irdy),
      .ivld(render_params_out_rsci_ivld_run_sct),
      .idat(render_params_out_rsci_idat),
      .rdy(render_params_out_rsc_rdy),
      .vld(render_params_out_rsc_vld),
      .dat(render_params_out_rsc_dat)
    );
  RenderLooper_run_render_params_out_rsci_render_params_out_wait_ctrl RenderLooper_run_render_params_out_rsci_render_params_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .render_params_out_rsci_oswt(render_params_out_rsci_oswt),
      .render_params_out_rsci_irdy(render_params_out_rsci_irdy),
      .render_params_out_rsci_biwt(render_params_out_rsci_biwt),
      .render_params_out_rsci_bdwt(render_params_out_rsci_bdwt),
      .render_params_out_rsci_bcwt(render_params_out_rsci_bcwt),
      .render_params_out_rsci_ivld_run_sct(render_params_out_rsci_ivld_run_sct)
    );
  RenderLooper_run_render_params_out_rsci_render_params_out_wait_dp RenderLooper_run_render_params_out_rsci_render_params_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_out_rsci_oswt(render_params_out_rsci_oswt),
      .render_params_out_rsci_wen_comp(render_params_out_rsci_wen_comp),
      .render_params_out_rsci_biwt(render_params_out_rsci_biwt),
      .render_params_out_rsci_bdwt(render_params_out_rsci_bdwt),
      .render_params_out_rsci_bcwt(render_params_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run_render_params_rsci
// ------------------------------------------------------------------


module RenderLooper_run_render_params_rsci (
  clk, arst_n, render_params_rsc_dat, render_params_rsc_vld, render_params_rsc_rdy,
      run_wen, render_params_rsci_oswt, render_params_rsci_wen_comp, render_params_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [419:0] render_params_rsc_dat;
  input render_params_rsc_vld;
  output render_params_rsc_rdy;
  input run_wen;
  input render_params_rsci_oswt;
  output render_params_rsci_wen_comp;
  output [419:0] render_params_rsci_idat_mxwt;


  // Interconnect Declarations
  wire render_params_rsci_biwt;
  wire render_params_rsci_bdwt;
  wire render_params_rsci_bcwt;
  wire render_params_rsci_irdy_run_sct;
  wire render_params_rsci_ivld;
  wire [419:0] render_params_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd21),
  .width(32'sd420)) render_params_rsci (
      .rdy(render_params_rsc_rdy),
      .vld(render_params_rsc_vld),
      .dat(render_params_rsc_dat),
      .irdy(render_params_rsci_irdy_run_sct),
      .ivld(render_params_rsci_ivld),
      .idat(render_params_rsci_idat)
    );
  RenderLooper_run_render_params_rsci_render_params_wait_ctrl RenderLooper_run_render_params_rsci_render_params_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .render_params_rsci_oswt(render_params_rsci_oswt),
      .render_params_rsci_biwt(render_params_rsci_biwt),
      .render_params_rsci_bdwt(render_params_rsci_bdwt),
      .render_params_rsci_bcwt(render_params_rsci_bcwt),
      .render_params_rsci_irdy_run_sct(render_params_rsci_irdy_run_sct),
      .render_params_rsci_ivld(render_params_rsci_ivld)
    );
  RenderLooper_run_render_params_rsci_render_params_wait_dp RenderLooper_run_render_params_rsci_render_params_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsci_oswt(render_params_rsci_oswt),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .render_params_rsci_idat_mxwt(render_params_rsci_idat_mxwt),
      .render_params_rsci_biwt(render_params_rsci_biwt),
      .render_params_rsci_bdwt(render_params_rsci_bdwt),
      .render_params_rsci_bcwt(render_params_rsci_bcwt),
      .render_params_rsci_idat(render_params_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_rayOut_rsci
// ------------------------------------------------------------------


module RayGeneration_run_rayOut_rsci (
  clk, arst_n, rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy, run_wen, rayOut_rsci_oswt,
      rayOut_rsci_wen_comp, rayOut_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;
  input run_wen;
  input rayOut_rsci_oswt;
  output rayOut_rsci_wen_comp;
  input [165:0] rayOut_rsci_idat;


  // Interconnect Declarations
  wire rayOut_rsci_irdy;
  wire rayOut_rsci_biwt;
  wire rayOut_rsci_bdwt;
  wire rayOut_rsci_bcwt;
  wire rayOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [165:0] nl_rayOut_rsci_idat;
  assign nl_rayOut_rsci_idat = {1'b1 , (rayOut_rsci_idat[164:132]) , 1'b0 , (rayOut_rsci_idat[130:98])
      , 1'b0 , (rayOut_rsci_idat[96:64]) , 1'b0 , (rayOut_rsci_idat[62:52]) , 10'b0000000000
      , (rayOut_rsci_idat[41:31]) , 10'b0000000000 , (rayOut_rsci_idat[20:10]) ,
      10'b0000000000};
  ccs_out_wait_v1 #(.rscid(32'sd27),
  .width(32'sd166)) rayOut_rsci (
      .irdy(rayOut_rsci_irdy),
      .ivld(rayOut_rsci_ivld_run_sct),
      .idat(nl_rayOut_rsci_idat[165:0]),
      .rdy(rayOut_rsc_rdy),
      .vld(rayOut_rsc_vld),
      .dat(rayOut_rsc_dat)
    );
  RayGeneration_run_rayOut_rsci_rayOut_wait_ctrl RayGeneration_run_rayOut_rsci_rayOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .rayOut_rsci_oswt(rayOut_rsci_oswt),
      .rayOut_rsci_irdy(rayOut_rsci_irdy),
      .rayOut_rsci_biwt(rayOut_rsci_biwt),
      .rayOut_rsci_bdwt(rayOut_rsci_bdwt),
      .rayOut_rsci_bcwt(rayOut_rsci_bcwt),
      .rayOut_rsci_ivld_run_sct(rayOut_rsci_ivld_run_sct)
    );
  RayGeneration_run_rayOut_rsci_rayOut_wait_dp RayGeneration_run_rayOut_rsci_rayOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rayOut_rsci_oswt(rayOut_rsci_oswt),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp),
      .rayOut_rsci_biwt(rayOut_rsci_biwt),
      .rayOut_rsci_bdwt(rayOut_rsci_bdwt),
      .rayOut_rsci_bcwt(rayOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsOut_rsci
// ------------------------------------------------------------------


module RayGeneration_run_paramsOut_rsci (
  clk, arst_n, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy, run_wen,
      paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_idat
);
  input clk;
  input arst_n;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  input run_wen;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input [92:0] paramsOut_rsci_idat;


  // Interconnect Declarations
  wire paramsOut_rsci_irdy;
  wire paramsOut_rsci_biwt;
  wire paramsOut_rsci_bdwt;
  wire paramsOut_rsci_bcwt;
  wire paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd26),
  .width(32'sd93)) paramsOut_rsci (
      .irdy(paramsOut_rsci_irdy),
      .ivld(paramsOut_rsci_ivld_run_sct),
      .idat(paramsOut_rsci_idat),
      .rdy(paramsOut_rsc_rdy),
      .vld(paramsOut_rsc_vld),
      .dat(paramsOut_rsc_dat)
    );
  RayGeneration_run_paramsOut_rsci_paramsOut_wait_ctrl RayGeneration_run_paramsOut_rsci_paramsOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_irdy(paramsOut_rsci_irdy),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt),
      .paramsOut_rsci_ivld_run_sct(paramsOut_rsci_ivld_run_sct)
    );
  RayGeneration_run_paramsOut_rsci_paramsOut_wait_dp RayGeneration_run_paramsOut_rsci_paramsOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_paramsIn_rsci
// ------------------------------------------------------------------


module RayGeneration_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [419:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [373:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [419:0] paramsIn_rsci_idat;
  wire [373:0] paramsIn_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd25),
  .width(32'sd420)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  RayGeneration_run_paramsIn_rsci_paramsIn_wait_ctrl RayGeneration_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  RayGeneration_run_paramsIn_rsci_paramsIn_wait_dp RayGeneration_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt_pconst),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
  assign paramsIn_rsci_idat_mxwt = paramsIn_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run_loopIndicesIn_rsci
// ------------------------------------------------------------------


module RayGeneration_run_loopIndicesIn_rsci (
  clk, arst_n, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld, loopIndicesIn_rsc_rdy,
      run_wen, loopIndicesIn_rsci_oswt, loopIndicesIn_rsci_wen_comp, loopIndicesIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [22:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  input run_wen;
  input loopIndicesIn_rsci_oswt;
  output loopIndicesIn_rsci_wen_comp;
  output [22:0] loopIndicesIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire loopIndicesIn_rsci_biwt;
  wire loopIndicesIn_rsci_bdwt;
  wire loopIndicesIn_rsci_bcwt;
  wire loopIndicesIn_rsci_irdy_run_sct;
  wire loopIndicesIn_rsci_ivld;
  wire [22:0] loopIndicesIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd24),
  .width(32'sd23)) loopIndicesIn_rsci (
      .rdy(loopIndicesIn_rsc_rdy),
      .vld(loopIndicesIn_rsc_vld),
      .dat(loopIndicesIn_rsc_dat),
      .irdy(loopIndicesIn_rsci_irdy_run_sct),
      .ivld(loopIndicesIn_rsci_ivld),
      .idat(loopIndicesIn_rsci_idat)
    );
  RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_irdy_run_sct(loopIndicesIn_rsci_irdy_run_sct),
      .loopIndicesIn_rsci_ivld(loopIndicesIn_rsci_ivld)
    );
  RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp RayGeneration_run_loopIndicesIn_rsci_loopIndicesIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsci_oswt(loopIndicesIn_rsci_oswt),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt),
      .loopIndicesIn_rsci_biwt(loopIndicesIn_rsci_biwt),
      .loopIndicesIn_rsci_bdwt(loopIndicesIn_rsci_bdwt),
      .loopIndicesIn_rsci_bcwt(loopIndicesIn_rsci_bcwt),
      .loopIndicesIn_rsci_idat(loopIndicesIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_out_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_params_out_rsci (
  clk, arst_n, params_out_rsc_dat, params_out_rsc_vld, params_out_rsc_rdy, run_wen,
      params_out_rsci_oswt, params_out_rsci_wen_comp, params_out_rsci_idat
);
  input clk;
  input arst_n;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;
  input run_wen;
  input params_out_rsci_oswt;
  output params_out_rsci_wen_comp;
  input [92:0] params_out_rsci_idat;


  // Interconnect Declarations
  wire params_out_rsci_irdy;
  wire params_out_rsci_biwt;
  wire params_out_rsci_bdwt;
  wire params_out_rsci_bcwt;
  wire params_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd42),
  .width(32'sd93)) params_out_rsci (
      .irdy(params_out_rsci_irdy),
      .ivld(params_out_rsci_ivld_run_sct),
      .idat(params_out_rsci_idat),
      .rdy(params_out_rsc_rdy),
      .vld(params_out_rsc_vld),
      .dat(params_out_rsc_dat)
    );
  LoopDistrib_run_params_out_rsci_params_out_wait_ctrl LoopDistrib_run_params_out_rsci_params_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .params_out_rsci_oswt(params_out_rsci_oswt),
      .params_out_rsci_irdy(params_out_rsci_irdy),
      .params_out_rsci_biwt(params_out_rsci_biwt),
      .params_out_rsci_bdwt(params_out_rsci_bdwt),
      .params_out_rsci_bcwt(params_out_rsci_bcwt),
      .params_out_rsci_ivld_run_sct(params_out_rsci_ivld_run_sct)
    );
  LoopDistrib_run_params_out_rsci_params_out_wait_dp LoopDistrib_run_params_out_rsci_params_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_out_rsci_oswt(params_out_rsci_oswt),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp),
      .params_out_rsci_biwt(params_out_rsci_biwt),
      .params_out_rsci_bdwt(params_out_rsci_bdwt),
      .params_out_rsci_bcwt(params_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outtwo_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outtwo_rsci (
  clk, arst_n, quad_max_outtwo_rsc_dat, quad_max_outtwo_rsc_vld, quad_max_outtwo_rsc_rdy,
      run_wen, quad_max_outtwo_rsci_oswt, quad_max_outtwo_rsci_wen_comp, quad_max_outtwo_rsci_idat
);
  input clk;
  input arst_n;
  output [10:0] quad_max_outtwo_rsc_dat;
  output quad_max_outtwo_rsc_vld;
  input quad_max_outtwo_rsc_rdy;
  input run_wen;
  input quad_max_outtwo_rsci_oswt;
  output quad_max_outtwo_rsci_wen_comp;
  input [10:0] quad_max_outtwo_rsci_idat;


  // Interconnect Declarations
  wire quad_max_outtwo_rsci_irdy;
  wire quad_max_outtwo_rsci_biwt;
  wire quad_max_outtwo_rsci_bdwt;
  wire quad_max_outtwo_rsci_bcwt;
  wire quad_max_outtwo_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd41),
  .width(32'sd11)) quad_max_outtwo_rsci (
      .irdy(quad_max_outtwo_rsci_irdy),
      .ivld(quad_max_outtwo_rsci_ivld_run_sct),
      .idat(quad_max_outtwo_rsci_idat),
      .rdy(quad_max_outtwo_rsc_rdy),
      .vld(quad_max_outtwo_rsc_vld),
      .dat(quad_max_outtwo_rsc_dat)
    );
  LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_ctrl LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quad_max_outtwo_rsci_oswt(quad_max_outtwo_rsci_oswt),
      .quad_max_outtwo_rsci_irdy(quad_max_outtwo_rsci_irdy),
      .quad_max_outtwo_rsci_biwt(quad_max_outtwo_rsci_biwt),
      .quad_max_outtwo_rsci_bdwt(quad_max_outtwo_rsci_bdwt),
      .quad_max_outtwo_rsci_bcwt(quad_max_outtwo_rsci_bcwt),
      .quad_max_outtwo_rsci_ivld_run_sct(quad_max_outtwo_rsci_ivld_run_sct)
    );
  LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_dp LoopDistrib_run_quad_max_outtwo_rsci_quad_max_outtwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_outtwo_rsci_oswt(quad_max_outtwo_rsci_oswt),
      .quad_max_outtwo_rsci_wen_comp(quad_max_outtwo_rsci_wen_comp),
      .quad_max_outtwo_rsci_biwt(quad_max_outtwo_rsci_biwt),
      .quad_max_outtwo_rsci_bdwt(quad_max_outtwo_rsci_bdwt),
      .quad_max_outtwo_rsci_bcwt(quad_max_outtwo_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_max_outone_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_quad_max_outone_rsci (
  clk, arst_n, quad_max_outone_rsc_dat, quad_max_outone_rsc_vld, quad_max_outone_rsc_rdy,
      run_wen, quad_max_outone_rsci_oswt, quad_max_outone_rsci_wen_comp, quad_max_outone_rsci_idat
);
  input clk;
  input arst_n;
  output [10:0] quad_max_outone_rsc_dat;
  output quad_max_outone_rsc_vld;
  input quad_max_outone_rsc_rdy;
  input run_wen;
  input quad_max_outone_rsci_oswt;
  output quad_max_outone_rsci_wen_comp;
  input [10:0] quad_max_outone_rsci_idat;


  // Interconnect Declarations
  wire quad_max_outone_rsci_irdy;
  wire quad_max_outone_rsci_biwt;
  wire quad_max_outone_rsci_bdwt;
  wire quad_max_outone_rsci_bcwt;
  wire quad_max_outone_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_quad_max_outone_rsci_idat;
  assign nl_quad_max_outone_rsci_idat = {1'b0 , (quad_max_outone_rsci_idat[9:0])};
  ccs_out_wait_v1 #(.rscid(32'sd40),
  .width(32'sd11)) quad_max_outone_rsci (
      .irdy(quad_max_outone_rsci_irdy),
      .ivld(quad_max_outone_rsci_ivld_run_sct),
      .idat(nl_quad_max_outone_rsci_idat[10:0]),
      .rdy(quad_max_outone_rsc_rdy),
      .vld(quad_max_outone_rsc_vld),
      .dat(quad_max_outone_rsc_dat)
    );
  LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_ctrl LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quad_max_outone_rsci_oswt(quad_max_outone_rsci_oswt),
      .quad_max_outone_rsci_irdy(quad_max_outone_rsci_irdy),
      .quad_max_outone_rsci_biwt(quad_max_outone_rsci_biwt),
      .quad_max_outone_rsci_bdwt(quad_max_outone_rsci_bdwt),
      .quad_max_outone_rsci_bcwt(quad_max_outone_rsci_bcwt),
      .quad_max_outone_rsci_ivld_run_sct(quad_max_outone_rsci_ivld_run_sct)
    );
  LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_dp LoopDistrib_run_quad_max_outone_rsci_quad_max_outone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_outone_rsci_oswt(quad_max_outone_rsci_oswt),
      .quad_max_outone_rsci_wen_comp(quad_max_outone_rsci_wen_comp),
      .quad_max_outone_rsci_biwt(quad_max_outone_rsci_biwt),
      .quad_max_outone_rsci_bdwt(quad_max_outone_rsci_bdwt),
      .quad_max_outone_rsci_bcwt(quad_max_outone_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_looptwo_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_looptwo_rsci (
  clk, arst_n, quad_out_looptwo_rsc_dat, quad_out_looptwo_rsc_vld, quad_out_looptwo_rsc_rdy,
      run_wen, quad_out_looptwo_rsci_oswt, quad_out_looptwo_rsci_wen_comp, quad_out_looptwo_rsci_idat
);
  input clk;
  input arst_n;
  output [376:0] quad_out_looptwo_rsc_dat;
  output quad_out_looptwo_rsc_vld;
  input quad_out_looptwo_rsc_rdy;
  input run_wen;
  input quad_out_looptwo_rsci_oswt;
  output quad_out_looptwo_rsci_wen_comp;
  input [376:0] quad_out_looptwo_rsci_idat;


  // Interconnect Declarations
  wire quad_out_looptwo_rsci_irdy;
  wire quad_out_looptwo_rsci_biwt;
  wire quad_out_looptwo_rsci_bdwt;
  wire quad_out_looptwo_rsci_bcwt;
  wire quad_out_looptwo_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd39),
  .width(32'sd377)) quad_out_looptwo_rsci (
      .irdy(quad_out_looptwo_rsci_irdy),
      .ivld(quad_out_looptwo_rsci_ivld_run_sct),
      .idat(quad_out_looptwo_rsci_idat),
      .rdy(quad_out_looptwo_rsc_rdy),
      .vld(quad_out_looptwo_rsc_vld),
      .dat(quad_out_looptwo_rsc_dat)
    );
  LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_ctrl LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quad_out_looptwo_rsci_oswt(quad_out_looptwo_rsci_oswt),
      .quad_out_looptwo_rsci_irdy(quad_out_looptwo_rsci_irdy),
      .quad_out_looptwo_rsci_biwt(quad_out_looptwo_rsci_biwt),
      .quad_out_looptwo_rsci_bdwt(quad_out_looptwo_rsci_bdwt),
      .quad_out_looptwo_rsci_bcwt(quad_out_looptwo_rsci_bcwt),
      .quad_out_looptwo_rsci_ivld_run_sct(quad_out_looptwo_rsci_ivld_run_sct)
    );
  LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_dp LoopDistrib_run_quad_out_looptwo_rsci_quad_out_looptwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_out_looptwo_rsci_oswt(quad_out_looptwo_rsci_oswt),
      .quad_out_looptwo_rsci_wen_comp(quad_out_looptwo_rsci_wen_comp),
      .quad_out_looptwo_rsci_biwt(quad_out_looptwo_rsci_biwt),
      .quad_out_looptwo_rsci_bdwt(quad_out_looptwo_rsci_bdwt),
      .quad_out_looptwo_rsci_bcwt(quad_out_looptwo_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quad_out_loopone_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_quad_out_loopone_rsci (
  clk, arst_n, quad_out_loopone_rsc_dat, quad_out_loopone_rsc_vld, quad_out_loopone_rsc_rdy,
      run_wen, quad_out_loopone_rsci_oswt, quad_out_loopone_rsci_wen_comp, quad_out_loopone_rsci_idat
);
  input clk;
  input arst_n;
  output [376:0] quad_out_loopone_rsc_dat;
  output quad_out_loopone_rsc_vld;
  input quad_out_loopone_rsc_rdy;
  input run_wen;
  input quad_out_loopone_rsci_oswt;
  output quad_out_loopone_rsci_wen_comp;
  input [376:0] quad_out_loopone_rsci_idat;


  // Interconnect Declarations
  wire quad_out_loopone_rsci_irdy;
  wire quad_out_loopone_rsci_biwt;
  wire quad_out_loopone_rsci_bdwt;
  wire quad_out_loopone_rsci_bcwt;
  wire quad_out_loopone_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd38),
  .width(32'sd377)) quad_out_loopone_rsci (
      .irdy(quad_out_loopone_rsci_irdy),
      .ivld(quad_out_loopone_rsci_ivld_run_sct),
      .idat(quad_out_loopone_rsci_idat),
      .rdy(quad_out_loopone_rsc_rdy),
      .vld(quad_out_loopone_rsc_vld),
      .dat(quad_out_loopone_rsc_dat)
    );
  LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_ctrl LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quad_out_loopone_rsci_oswt(quad_out_loopone_rsci_oswt),
      .quad_out_loopone_rsci_irdy(quad_out_loopone_rsci_irdy),
      .quad_out_loopone_rsci_biwt(quad_out_loopone_rsci_biwt),
      .quad_out_loopone_rsci_bdwt(quad_out_loopone_rsci_bdwt),
      .quad_out_loopone_rsci_bcwt(quad_out_loopone_rsci_bcwt),
      .quad_out_loopone_rsci_ivld_run_sct(quad_out_loopone_rsci_ivld_run_sct)
    );
  LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_dp LoopDistrib_run_quad_out_loopone_rsci_quad_out_loopone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_out_loopone_rsci_oswt(quad_out_loopone_rsci_oswt),
      .quad_out_loopone_rsci_wen_comp(quad_out_loopone_rsci_wen_comp),
      .quad_out_loopone_rsci_biwt(quad_out_loopone_rsci_biwt),
      .quad_out_loopone_rsci_bdwt(quad_out_loopone_rsci_bdwt),
      .quad_out_loopone_rsci_bcwt(quad_out_loopone_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_worldhit_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_worldhit_rsci (
  clk, arst_n, ray_out_worldhit_rsc_dat, ray_out_worldhit_rsc_vld, ray_out_worldhit_rsc_rdy,
      run_wen, ray_out_worldhit_rsci_oswt, ray_out_worldhit_rsci_wen_comp, ray_out_worldhit_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_worldhit_rsc_dat;
  output ray_out_worldhit_rsc_vld;
  input ray_out_worldhit_rsc_rdy;
  input run_wen;
  input ray_out_worldhit_rsci_oswt;
  output ray_out_worldhit_rsci_wen_comp;
  input [165:0] ray_out_worldhit_rsci_idat;


  // Interconnect Declarations
  wire ray_out_worldhit_rsci_irdy;
  wire ray_out_worldhit_rsci_biwt;
  wire ray_out_worldhit_rsci_bdwt;
  wire ray_out_worldhit_rsci_bcwt;
  wire ray_out_worldhit_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd37),
  .width(32'sd166)) ray_out_worldhit_rsci (
      .irdy(ray_out_worldhit_rsci_irdy),
      .ivld(ray_out_worldhit_rsci_ivld_run_sct),
      .idat(ray_out_worldhit_rsci_idat),
      .rdy(ray_out_worldhit_rsc_rdy),
      .vld(ray_out_worldhit_rsc_vld),
      .dat(ray_out_worldhit_rsc_dat)
    );
  LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_ctrl LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_out_worldhit_rsci_oswt(ray_out_worldhit_rsci_oswt),
      .ray_out_worldhit_rsci_irdy(ray_out_worldhit_rsci_irdy),
      .ray_out_worldhit_rsci_biwt(ray_out_worldhit_rsci_biwt),
      .ray_out_worldhit_rsci_bdwt(ray_out_worldhit_rsci_bdwt),
      .ray_out_worldhit_rsci_bcwt(ray_out_worldhit_rsci_bcwt),
      .ray_out_worldhit_rsci_ivld_run_sct(ray_out_worldhit_rsci_ivld_run_sct)
    );
  LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_dp LoopDistrib_run_ray_out_worldhit_rsci_ray_out_worldhit_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_worldhit_rsci_oswt(ray_out_worldhit_rsci_oswt),
      .ray_out_worldhit_rsci_wen_comp(ray_out_worldhit_rsci_wen_comp),
      .ray_out_worldhit_rsci_biwt(ray_out_worldhit_rsci_biwt),
      .ray_out_worldhit_rsci_bdwt(ray_out_worldhit_rsci_bdwt),
      .ray_out_worldhit_rsci_bcwt(ray_out_worldhit_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_looptwo_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_looptwo_rsci (
  clk, arst_n, ray_out_looptwo_rsc_dat, ray_out_looptwo_rsc_vld, ray_out_looptwo_rsc_rdy,
      run_wen, ray_out_looptwo_rsci_oswt, ray_out_looptwo_rsci_wen_comp, ray_out_looptwo_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_looptwo_rsc_dat;
  output ray_out_looptwo_rsc_vld;
  input ray_out_looptwo_rsc_rdy;
  input run_wen;
  input ray_out_looptwo_rsci_oswt;
  output ray_out_looptwo_rsci_wen_comp;
  input [165:0] ray_out_looptwo_rsci_idat;


  // Interconnect Declarations
  wire ray_out_looptwo_rsci_irdy;
  wire ray_out_looptwo_rsci_biwt;
  wire ray_out_looptwo_rsci_bdwt;
  wire ray_out_looptwo_rsci_bcwt;
  wire ray_out_looptwo_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd36),
  .width(32'sd166)) ray_out_looptwo_rsci (
      .irdy(ray_out_looptwo_rsci_irdy),
      .ivld(ray_out_looptwo_rsci_ivld_run_sct),
      .idat(ray_out_looptwo_rsci_idat),
      .rdy(ray_out_looptwo_rsc_rdy),
      .vld(ray_out_looptwo_rsc_vld),
      .dat(ray_out_looptwo_rsc_dat)
    );
  LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_ctrl LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_out_looptwo_rsci_oswt(ray_out_looptwo_rsci_oswt),
      .ray_out_looptwo_rsci_irdy(ray_out_looptwo_rsci_irdy),
      .ray_out_looptwo_rsci_biwt(ray_out_looptwo_rsci_biwt),
      .ray_out_looptwo_rsci_bdwt(ray_out_looptwo_rsci_bdwt),
      .ray_out_looptwo_rsci_bcwt(ray_out_looptwo_rsci_bcwt),
      .ray_out_looptwo_rsci_ivld_run_sct(ray_out_looptwo_rsci_ivld_run_sct)
    );
  LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_dp LoopDistrib_run_ray_out_looptwo_rsci_ray_out_looptwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_looptwo_rsci_oswt(ray_out_looptwo_rsci_oswt),
      .ray_out_looptwo_rsci_wen_comp(ray_out_looptwo_rsci_wen_comp),
      .ray_out_looptwo_rsci_biwt(ray_out_looptwo_rsci_biwt),
      .ray_out_looptwo_rsci_bdwt(ray_out_looptwo_rsci_bdwt),
      .ray_out_looptwo_rsci_bcwt(ray_out_looptwo_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_out_loopone_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_ray_out_loopone_rsci (
  clk, arst_n, ray_out_loopone_rsc_dat, ray_out_loopone_rsc_vld, ray_out_loopone_rsc_rdy,
      run_wen, ray_out_loopone_rsci_oswt, ray_out_loopone_rsci_wen_comp, ray_out_loopone_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_loopone_rsc_dat;
  output ray_out_loopone_rsc_vld;
  input ray_out_loopone_rsc_rdy;
  input run_wen;
  input ray_out_loopone_rsci_oswt;
  output ray_out_loopone_rsci_wen_comp;
  input [165:0] ray_out_loopone_rsci_idat;


  // Interconnect Declarations
  wire ray_out_loopone_rsci_irdy;
  wire ray_out_loopone_rsci_biwt;
  wire ray_out_loopone_rsci_bdwt;
  wire ray_out_loopone_rsci_bcwt;
  wire ray_out_loopone_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd35),
  .width(32'sd166)) ray_out_loopone_rsci (
      .irdy(ray_out_loopone_rsci_irdy),
      .ivld(ray_out_loopone_rsci_ivld_run_sct),
      .idat(ray_out_loopone_rsci_idat),
      .rdy(ray_out_loopone_rsc_rdy),
      .vld(ray_out_loopone_rsc_vld),
      .dat(ray_out_loopone_rsc_dat)
    );
  LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_ctrl LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_out_loopone_rsci_oswt(ray_out_loopone_rsci_oswt),
      .ray_out_loopone_rsci_irdy(ray_out_loopone_rsci_irdy),
      .ray_out_loopone_rsci_biwt(ray_out_loopone_rsci_biwt),
      .ray_out_loopone_rsci_bdwt(ray_out_loopone_rsci_bdwt),
      .ray_out_loopone_rsci_bcwt(ray_out_loopone_rsci_bcwt),
      .ray_out_loopone_rsci_ivld_run_sct(ray_out_loopone_rsci_ivld_run_sct)
    );
  LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_dp LoopDistrib_run_ray_out_loopone_rsci_ray_out_loopone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_loopone_rsci_oswt(ray_out_loopone_rsci_oswt),
      .ray_out_loopone_rsci_wen_comp(ray_out_loopone_rsci_wen_comp),
      .ray_out_loopone_rsci_biwt(ray_out_loopone_rsci_biwt),
      .ray_out_loopone_rsci_bdwt(ray_out_loopone_rsci_bdwt),
      .ray_out_loopone_rsci_bcwt(ray_out_loopone_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_out_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_out_rsci (
  clk, arst_n, accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      run_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  input run_wen;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input [80:0] accumalated_color_out_rsci_idat;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_irdy;
  wire accumalated_color_out_rsci_biwt;
  wire accumalated_color_out_rsci_bdwt;
  wire accumalated_color_out_rsci_bcwt;
  wire accumalated_color_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd34),
  .width(32'sd81)) accumalated_color_out_rsci (
      .irdy(accumalated_color_out_rsci_irdy),
      .ivld(accumalated_color_out_rsci_ivld_run_sct),
      .idat(accumalated_color_out_rsci_idat),
      .rdy(accumalated_color_out_rsc_rdy),
      .vld(accumalated_color_out_rsc_vld),
      .dat(accumalated_color_out_rsc_dat)
    );
  LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_irdy(accumalated_color_out_rsci_irdy),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt),
      .accumalated_color_out_rsci_ivld_run_sct(accumalated_color_out_rsci_ivld_run_sct)
    );
  LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_dp LoopDistrib_run_accumalated_color_out_rsci_accumalated_color_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_out_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_out_rsci (
  clk, arst_n, attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      run_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  input run_wen;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input [80:0] attenuation_chan_out_rsci_idat;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_irdy;
  wire attenuation_chan_out_rsci_biwt;
  wire attenuation_chan_out_rsci_bdwt;
  wire attenuation_chan_out_rsci_bcwt;
  wire attenuation_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd33),
  .width(32'sd81)) attenuation_chan_out_rsci (
      .irdy(attenuation_chan_out_rsci_irdy),
      .ivld(attenuation_chan_out_rsci_ivld_run_sct),
      .idat(attenuation_chan_out_rsci_idat),
      .rdy(attenuation_chan_out_rsc_rdy),
      .vld(attenuation_chan_out_rsc_vld),
      .dat(attenuation_chan_out_rsc_dat)
    );
  LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_irdy(attenuation_chan_out_rsci_irdy),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt),
      .attenuation_chan_out_rsci_ivld_run_sct(attenuation_chan_out_rsci_ivld_run_sct)
    );
  LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp LoopDistrib_run_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_accumalated_color_chan_in_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_accumalated_color_chan_in_rsci (
  clk, arst_n, accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld,
      accumalated_color_chan_in_rsc_rdy, run_wen, accumalated_color_chan_in_rsci_oswt,
      accumalated_color_chan_in_rsci_wen_comp, accumalated_color_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input run_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_biwt;
  wire accumalated_color_chan_in_rsci_bdwt;
  wire accumalated_color_chan_in_rsci_bcwt;
  wire accumalated_color_chan_in_rsci_irdy_run_sct;
  wire accumalated_color_chan_in_rsci_ivld;
  wire [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd32),
  .width(32'sd81)) accumalated_color_chan_in_rsci (
      .rdy(accumalated_color_chan_in_rsc_rdy),
      .vld(accumalated_color_chan_in_rsc_vld),
      .dat(accumalated_color_chan_in_rsc_dat),
      .irdy(accumalated_color_chan_in_rsci_irdy_run_sct),
      .ivld(accumalated_color_chan_in_rsci_ivld),
      .idat(accumalated_color_chan_in_rsci_idat)
    );
  LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
      LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_irdy_run_sct(accumalated_color_chan_in_rsci_irdy_run_sct),
      .accumalated_color_chan_in_rsci_ivld(accumalated_color_chan_in_rsci_ivld)
    );
  LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
      LoopDistrib_run_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_idat(accumalated_color_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_attenuation_chan_in_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_attenuation_chan_in_rsci (
  clk, arst_n, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      run_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input run_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_biwt;
  wire attenuation_chan_in_rsci_bdwt;
  wire attenuation_chan_in_rsci_bcwt;
  wire attenuation_chan_in_rsci_irdy_run_sct;
  wire attenuation_chan_in_rsci_ivld;
  wire [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd31),
  .width(32'sd81)) attenuation_chan_in_rsci (
      .rdy(attenuation_chan_in_rsc_rdy),
      .vld(attenuation_chan_in_rsc_vld),
      .dat(attenuation_chan_in_rsc_dat),
      .irdy(attenuation_chan_in_rsci_irdy_run_sct),
      .ivld(attenuation_chan_in_rsci_ivld),
      .idat(attenuation_chan_in_rsci_idat)
    );
  LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_irdy_run_sct(attenuation_chan_in_rsci_irdy_run_sct),
      .attenuation_chan_in_rsci_ivld(attenuation_chan_in_rsci_ivld)
    );
  LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp LoopDistrib_run_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_idat(attenuation_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_quads_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_quads_rsci (
  clk, arst_n, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy, run_wen, quads_rsci_oswt,
      quads_rsci_wen_comp, quads_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input run_wen;
  input quads_rsci_oswt;
  output quads_rsci_wen_comp;
  output [376:0] quads_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quads_rsci_biwt;
  wire quads_rsci_bdwt;
  wire quads_rsci_bcwt;
  wire quads_rsci_irdy_run_sct;
  wire quads_rsci_ivld;
  wire [376:0] quads_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd30),
  .width(32'sd377)) quads_rsci (
      .rdy(quads_rsc_rdy),
      .vld(quads_rsc_vld),
      .dat(quads_rsc_dat),
      .irdy(quads_rsci_irdy_run_sct),
      .ivld(quads_rsci_ivld),
      .idat(quads_rsci_idat)
    );
  LoopDistrib_run_quads_rsci_quads_wait_ctrl LoopDistrib_run_quads_rsci_quads_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .quads_rsci_oswt(quads_rsci_oswt),
      .quads_rsci_biwt(quads_rsci_biwt),
      .quads_rsci_bdwt(quads_rsci_bdwt),
      .quads_rsci_bcwt(quads_rsci_bcwt),
      .quads_rsci_irdy_run_sct(quads_rsci_irdy_run_sct),
      .quads_rsci_ivld(quads_rsci_ivld)
    );
  LoopDistrib_run_quads_rsci_quads_wait_dp LoopDistrib_run_quads_rsci_quads_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsci_oswt(quads_rsci_oswt),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .quads_rsci_idat_mxwt(quads_rsci_idat_mxwt),
      .quads_rsci_biwt(quads_rsci_biwt),
      .quads_rsci_bdwt(quads_rsci_bdwt),
      .quads_rsci_bcwt(quads_rsci_bcwt),
      .quads_rsci_idat(quads_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_params_in_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_params_in_rsci (
  clk, arst_n, params_in_rsc_dat, params_in_rsc_vld, params_in_rsc_rdy, run_wen,
      params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input run_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [92:0] params_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire params_in_rsci_biwt;
  wire params_in_rsci_bdwt;
  wire params_in_rsci_bcwt;
  wire params_in_rsci_irdy_run_sct;
  wire params_in_rsci_ivld;
  wire [92:0] params_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd29),
  .width(32'sd93)) params_in_rsci (
      .rdy(params_in_rsc_rdy),
      .vld(params_in_rsc_vld),
      .dat(params_in_rsc_dat),
      .irdy(params_in_rsci_irdy_run_sct),
      .ivld(params_in_rsci_ivld),
      .idat(params_in_rsci_idat)
    );
  LoopDistrib_run_params_in_rsci_params_in_wait_ctrl LoopDistrib_run_params_in_rsci_params_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_irdy_run_sct(params_in_rsci_irdy_run_sct),
      .params_in_rsci_ivld(params_in_rsci_ivld)
    );
  LoopDistrib_run_params_in_rsci_params_in_wait_dp LoopDistrib_run_params_in_rsci_params_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_idat(params_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run_ray_in_rsci
// ------------------------------------------------------------------


module LoopDistrib_run_ray_in_rsci (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, run_wen, ray_in_rsci_oswt,
      ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input run_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [165:0] ray_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_in_rsci_biwt;
  wire ray_in_rsci_bdwt;
  wire ray_in_rsci_bcwt;
  wire ray_in_rsci_irdy_run_sct;
  wire ray_in_rsci_ivld;
  wire [165:0] ray_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd28),
  .width(32'sd166)) ray_in_rsci (
      .rdy(ray_in_rsc_rdy),
      .vld(ray_in_rsc_vld),
      .dat(ray_in_rsc_dat),
      .irdy(ray_in_rsci_irdy_run_sct),
      .ivld(ray_in_rsci_ivld),
      .idat(ray_in_rsci_idat)
    );
  LoopDistrib_run_ray_in_rsci_ray_in_wait_ctrl LoopDistrib_run_ray_in_rsci_ray_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_irdy_run_sct(ray_in_rsci_irdy_run_sct),
      .ray_in_rsci_ivld(ray_in_rsci_ivld)
    );
  LoopDistrib_run_ray_in_rsci_ray_in_wait_dp LoopDistrib_run_ray_in_rsci_ray_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_idat(ray_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_closest_so_far_out_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_closest_so_far_out_rsci (
  clk, arst_n, closest_so_far_out_rsc_dat, closest_so_far_out_rsc_vld, closest_so_far_out_rsc_rdy,
      hit_wen, closest_so_far_out_rsci_oswt, closest_so_far_out_rsci_wen_comp, closest_so_far_out_rsci_idat
);
  input clk;
  input arst_n;
  output [46:0] closest_so_far_out_rsc_dat;
  output closest_so_far_out_rsc_vld;
  input closest_so_far_out_rsc_rdy;
  input hit_wen;
  input closest_so_far_out_rsci_oswt;
  output closest_so_far_out_rsci_wen_comp;
  input [46:0] closest_so_far_out_rsci_idat;


  // Interconnect Declarations
  wire closest_so_far_out_rsci_irdy;
  wire closest_so_far_out_rsci_biwt;
  wire closest_so_far_out_rsci_bdwt;
  wire closest_so_far_out_rsci_bcwt;
  wire closest_so_far_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd48),
  .width(32'sd47)) closest_so_far_out_rsci (
      .irdy(closest_so_far_out_rsci_irdy),
      .ivld(closest_so_far_out_rsci_ivld_hit_sct),
      .idat(closest_so_far_out_rsci_idat),
      .rdy(closest_so_far_out_rsc_rdy),
      .vld(closest_so_far_out_rsc_vld),
      .dat(closest_so_far_out_rsc_dat)
    );
  IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_ctrl IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .closest_so_far_out_rsci_oswt(closest_so_far_out_rsci_oswt),
      .closest_so_far_out_rsci_irdy(closest_so_far_out_rsci_irdy),
      .closest_so_far_out_rsci_biwt(closest_so_far_out_rsci_biwt),
      .closest_so_far_out_rsci_bdwt(closest_so_far_out_rsci_bdwt),
      .closest_so_far_out_rsci_bcwt(closest_so_far_out_rsci_bcwt),
      .closest_so_far_out_rsci_ivld_hit_sct(closest_so_far_out_rsci_ivld_hit_sct)
    );
  IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_dp IntersecLoop_hit_closest_so_far_out_rsci_closest_so_far_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_out_rsci_oswt(closest_so_far_out_rsci_oswt),
      .closest_so_far_out_rsci_wen_comp(closest_so_far_out_rsci_wen_comp),
      .closest_so_far_out_rsci_biwt(closest_so_far_out_rsci_biwt),
      .closest_so_far_out_rsci_bdwt(closest_so_far_out_rsci_bdwt),
      .closest_so_far_out_rsci_bcwt(closest_so_far_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_rec_quad_out_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_rec_quad_out_rsci (
  clk, arst_n, rec_quad_out_rsc_dat, rec_quad_out_rsc_vld, rec_quad_out_rsc_rdy,
      hit_wen, rec_quad_out_rsci_oswt, rec_quad_out_rsci_wen_comp, rec_quad_out_rsci_idat
);
  input clk;
  input arst_n;
  output [225:0] rec_quad_out_rsc_dat;
  output rec_quad_out_rsc_vld;
  input rec_quad_out_rsc_rdy;
  input hit_wen;
  input rec_quad_out_rsci_oswt;
  output rec_quad_out_rsci_wen_comp;
  input [225:0] rec_quad_out_rsci_idat;


  // Interconnect Declarations
  wire rec_quad_out_rsci_irdy;
  wire rec_quad_out_rsci_biwt;
  wire rec_quad_out_rsci_bdwt;
  wire rec_quad_out_rsci_bcwt;
  wire rec_quad_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd47),
  .width(32'sd226)) rec_quad_out_rsci (
      .irdy(rec_quad_out_rsci_irdy),
      .ivld(rec_quad_out_rsci_ivld_hit_sct),
      .idat(rec_quad_out_rsci_idat),
      .rdy(rec_quad_out_rsc_rdy),
      .vld(rec_quad_out_rsc_vld),
      .dat(rec_quad_out_rsc_dat)
    );
  IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_ctrl IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .rec_quad_out_rsci_oswt(rec_quad_out_rsci_oswt),
      .rec_quad_out_rsci_irdy(rec_quad_out_rsci_irdy),
      .rec_quad_out_rsci_biwt(rec_quad_out_rsci_biwt),
      .rec_quad_out_rsci_bdwt(rec_quad_out_rsci_bdwt),
      .rec_quad_out_rsci_bcwt(rec_quad_out_rsci_bcwt),
      .rec_quad_out_rsci_ivld_hit_sct(rec_quad_out_rsci_ivld_hit_sct)
    );
  IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_dp IntersecLoop_hit_rec_quad_out_rsci_rec_quad_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_out_rsci_oswt(rec_quad_out_rsci_oswt),
      .rec_quad_out_rsci_wen_comp(rec_quad_out_rsci_wen_comp),
      .rec_quad_out_rsci_biwt(rec_quad_out_rsci_biwt),
      .rec_quad_out_rsci_bdwt(rec_quad_out_rsci_bdwt),
      .rec_quad_out_rsci_bcwt(rec_quad_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_hit_anything_out_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_hit_anything_out_rsci (
  clk, arst_n, quad_hit_anything_out_rsc_dat, quad_hit_anything_out_rsc_vld, quad_hit_anything_out_rsc_rdy,
      hit_wen, quad_hit_anything_out_rsci_oswt, quad_hit_anything_out_rsci_wen_comp,
      quad_hit_anything_out_rsci_idat
);
  input clk;
  input arst_n;
  output quad_hit_anything_out_rsc_dat;
  output quad_hit_anything_out_rsc_vld;
  input quad_hit_anything_out_rsc_rdy;
  input hit_wen;
  input quad_hit_anything_out_rsci_oswt;
  output quad_hit_anything_out_rsci_wen_comp;
  input quad_hit_anything_out_rsci_idat;


  // Interconnect Declarations
  wire quad_hit_anything_out_rsci_irdy;
  wire quad_hit_anything_out_rsci_biwt;
  wire quad_hit_anything_out_rsci_bdwt;
  wire quad_hit_anything_out_rsci_bcwt;
  wire quad_hit_anything_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd46),
  .width(32'sd1)) quad_hit_anything_out_rsci (
      .irdy(quad_hit_anything_out_rsci_irdy),
      .ivld(quad_hit_anything_out_rsci_ivld_hit_sct),
      .idat(quad_hit_anything_out_rsci_idat),
      .rdy(quad_hit_anything_out_rsc_rdy),
      .vld(quad_hit_anything_out_rsc_vld),
      .dat(quad_hit_anything_out_rsc_dat)
    );
  IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_ctrl IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .quad_hit_anything_out_rsci_oswt(quad_hit_anything_out_rsci_oswt),
      .quad_hit_anything_out_rsci_irdy(quad_hit_anything_out_rsci_irdy),
      .quad_hit_anything_out_rsci_biwt(quad_hit_anything_out_rsci_biwt),
      .quad_hit_anything_out_rsci_bdwt(quad_hit_anything_out_rsci_bdwt),
      .quad_hit_anything_out_rsci_bcwt(quad_hit_anything_out_rsci_bcwt),
      .quad_hit_anything_out_rsci_ivld_hit_sct(quad_hit_anything_out_rsci_ivld_hit_sct)
    );
  IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_dp IntersecLoop_hit_quad_hit_anything_out_rsci_quad_hit_anything_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_out_rsci_oswt(quad_hit_anything_out_rsci_oswt),
      .quad_hit_anything_out_rsci_wen_comp(quad_hit_anything_out_rsci_wen_comp),
      .quad_hit_anything_out_rsci_biwt(quad_hit_anything_out_rsci_biwt),
      .quad_hit_anything_out_rsci_bdwt(quad_hit_anything_out_rsci_bdwt),
      .quad_hit_anything_out_rsci_bcwt(quad_hit_anything_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quad_max_in_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_quad_max_in_rsci (
  clk, arst_n, quad_max_in_rsc_dat, quad_max_in_rsc_vld, quad_max_in_rsc_rdy, hit_wen,
      quad_max_in_rsci_oswt, quad_max_in_rsci_wen_comp, quad_max_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [10:0] quad_max_in_rsc_dat;
  input quad_max_in_rsc_vld;
  output quad_max_in_rsc_rdy;
  input hit_wen;
  input quad_max_in_rsci_oswt;
  output quad_max_in_rsci_wen_comp;
  output [10:0] quad_max_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quad_max_in_rsci_biwt;
  wire quad_max_in_rsci_bdwt;
  wire quad_max_in_rsci_bcwt;
  wire quad_max_in_rsci_irdy_hit_sct;
  wire quad_max_in_rsci_ivld;
  wire [10:0] quad_max_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd45),
  .width(32'sd11)) quad_max_in_rsci (
      .rdy(quad_max_in_rsc_rdy),
      .vld(quad_max_in_rsc_vld),
      .dat(quad_max_in_rsc_dat),
      .irdy(quad_max_in_rsci_irdy_hit_sct),
      .ivld(quad_max_in_rsci_ivld),
      .idat(quad_max_in_rsci_idat)
    );
  IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_ctrl IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .quad_max_in_rsci_oswt(quad_max_in_rsci_oswt),
      .quad_max_in_rsci_biwt(quad_max_in_rsci_biwt),
      .quad_max_in_rsci_bdwt(quad_max_in_rsci_bdwt),
      .quad_max_in_rsci_bcwt(quad_max_in_rsci_bcwt),
      .quad_max_in_rsci_irdy_hit_sct(quad_max_in_rsci_irdy_hit_sct),
      .quad_max_in_rsci_ivld(quad_max_in_rsci_ivld)
    );
  IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_dp IntersecLoop_hit_quad_max_in_rsci_quad_max_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_in_rsci_oswt(quad_max_in_rsci_oswt),
      .quad_max_in_rsci_wen_comp(quad_max_in_rsci_wen_comp),
      .quad_max_in_rsci_idat_mxwt(quad_max_in_rsci_idat_mxwt),
      .quad_max_in_rsci_biwt(quad_max_in_rsci_biwt),
      .quad_max_in_rsci_bdwt(quad_max_in_rsci_bdwt),
      .quad_max_in_rsci_bcwt(quad_max_in_rsci_bcwt),
      .quad_max_in_rsci_idat(quad_max_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_ray_temp_in_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_ray_temp_in_rsci (
  clk, arst_n, ray_temp_in_rsc_dat, ray_temp_in_rsc_vld, ray_temp_in_rsc_rdy, hit_wen,
      ray_temp_in_rsci_oswt, ray_temp_in_rsci_wen_comp, ray_temp_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_temp_in_rsc_dat;
  input ray_temp_in_rsc_vld;
  output ray_temp_in_rsc_rdy;
  input hit_wen;
  input ray_temp_in_rsci_oswt;
  output ray_temp_in_rsci_wen_comp;
  output [165:0] ray_temp_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_temp_in_rsci_biwt;
  wire ray_temp_in_rsci_bdwt;
  wire ray_temp_in_rsci_bcwt;
  wire ray_temp_in_rsci_irdy_hit_sct;
  wire ray_temp_in_rsci_ivld;
  wire [165:0] ray_temp_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd44),
  .width(32'sd166)) ray_temp_in_rsci (
      .rdy(ray_temp_in_rsc_rdy),
      .vld(ray_temp_in_rsc_vld),
      .dat(ray_temp_in_rsc_dat),
      .irdy(ray_temp_in_rsci_irdy_hit_sct),
      .ivld(ray_temp_in_rsci_ivld),
      .idat(ray_temp_in_rsci_idat)
    );
  IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_ctrl IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .ray_temp_in_rsci_oswt(ray_temp_in_rsci_oswt),
      .ray_temp_in_rsci_biwt(ray_temp_in_rsci_biwt),
      .ray_temp_in_rsci_bdwt(ray_temp_in_rsci_bdwt),
      .ray_temp_in_rsci_bcwt(ray_temp_in_rsci_bcwt),
      .ray_temp_in_rsci_irdy_hit_sct(ray_temp_in_rsci_irdy_hit_sct),
      .ray_temp_in_rsci_ivld(ray_temp_in_rsci_ivld)
    );
  IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_dp IntersecLoop_hit_ray_temp_in_rsci_ray_temp_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_temp_in_rsci_oswt(ray_temp_in_rsci_oswt),
      .ray_temp_in_rsci_wen_comp(ray_temp_in_rsci_wen_comp),
      .ray_temp_in_rsci_idat_mxwt(ray_temp_in_rsci_idat_mxwt),
      .ray_temp_in_rsci_biwt(ray_temp_in_rsci_biwt),
      .ray_temp_in_rsci_bdwt(ray_temp_in_rsci_bdwt),
      .ray_temp_in_rsci_bcwt(ray_temp_in_rsci_bcwt),
      .ray_temp_in_rsci_idat(ray_temp_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit_quads_rsci
// ------------------------------------------------------------------


module IntersecLoop_hit_quads_rsci (
  clk, arst_n, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy, hit_wen, quads_rsci_oswt,
      quads_rsci_wen_comp, quads_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input hit_wen;
  input quads_rsci_oswt;
  output quads_rsci_wen_comp;
  output [376:0] quads_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quads_rsci_biwt;
  wire quads_rsci_bdwt;
  wire quads_rsci_bcwt;
  wire quads_rsci_irdy_hit_sct;
  wire quads_rsci_ivld;
  wire [376:0] quads_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd43),
  .width(32'sd377)) quads_rsci (
      .rdy(quads_rsc_rdy),
      .vld(quads_rsc_vld),
      .dat(quads_rsc_dat),
      .irdy(quads_rsci_irdy_hit_sct),
      .ivld(quads_rsci_ivld),
      .idat(quads_rsci_idat)
    );
  IntersecLoop_hit_quads_rsci_quads_wait_ctrl IntersecLoop_hit_quads_rsci_quads_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .quads_rsci_oswt(quads_rsci_oswt),
      .quads_rsci_biwt(quads_rsci_biwt),
      .quads_rsci_bdwt(quads_rsci_bdwt),
      .quads_rsci_bcwt(quads_rsci_bcwt),
      .quads_rsci_irdy_hit_sct(quads_rsci_irdy_hit_sct),
      .quads_rsci_ivld(quads_rsci_ivld)
    );
  IntersecLoop_hit_quads_rsci_quads_wait_dp IntersecLoop_hit_quads_rsci_quads_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsci_oswt(quads_rsci_oswt),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .quads_rsci_idat_mxwt(quads_rsci_idat_mxwt),
      .quads_rsci_biwt(quads_rsci_biwt),
      .quads_rsci_bdwt(quads_rsci_bdwt),
      .quads_rsci_bcwt(quads_rsci_bcwt),
      .quads_rsci_idat(quads_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_isHit_rsci
// ------------------------------------------------------------------


module WorldHit_hit_isHit_rsci (
  clk, arst_n, isHit_rsc_dat, isHit_rsc_vld, isHit_rsc_rdy, hit_wen, isHit_rsci_oswt,
      isHit_rsci_wen_comp, isHit_rsci_idat
);
  input clk;
  input arst_n;
  output isHit_rsc_dat;
  output isHit_rsc_vld;
  input isHit_rsc_rdy;
  input hit_wen;
  input isHit_rsci_oswt;
  output isHit_rsci_wen_comp;
  input isHit_rsci_idat;


  // Interconnect Declarations
  wire isHit_rsci_irdy;
  wire isHit_rsci_biwt;
  wire isHit_rsci_bdwt;
  wire isHit_rsci_bcwt;
  wire isHit_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd63),
  .width(32'sd1)) isHit_rsci (
      .irdy(isHit_rsci_irdy),
      .ivld(isHit_rsci_ivld_hit_sct),
      .idat(isHit_rsci_idat),
      .rdy(isHit_rsc_rdy),
      .vld(isHit_rsc_vld),
      .dat(isHit_rsc_dat)
    );
  WorldHit_hit_isHit_rsci_isHit_wait_ctrl WorldHit_hit_isHit_rsci_isHit_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .isHit_rsci_oswt(isHit_rsci_oswt),
      .isHit_rsci_irdy(isHit_rsci_irdy),
      .isHit_rsci_biwt(isHit_rsci_biwt),
      .isHit_rsci_bdwt(isHit_rsci_bdwt),
      .isHit_rsci_bcwt(isHit_rsci_bcwt),
      .isHit_rsci_ivld_hit_sct(isHit_rsci_ivld_hit_sct)
    );
  WorldHit_hit_isHit_rsci_isHit_wait_dp WorldHit_hit_isHit_rsci_isHit_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .isHit_rsci_oswt(isHit_rsci_oswt),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp),
      .isHit_rsci_biwt(isHit_rsci_biwt),
      .isHit_rsci_bdwt(isHit_rsci_bdwt),
      .isHit_rsci_bcwt(isHit_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_out_rsci
// ------------------------------------------------------------------


module WorldHit_hit_ray_out_rsci (
  clk, arst_n, ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, hit_wen, ray_out_rsci_oswt,
      ray_out_rsci_wen_comp, ray_out_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  input hit_wen;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input [165:0] ray_out_rsci_idat;


  // Interconnect Declarations
  wire ray_out_rsci_irdy;
  wire ray_out_rsci_biwt;
  wire ray_out_rsci_bdwt;
  wire ray_out_rsci_bcwt;
  wire ray_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  wire [165:0] nl_ray_out_rsci_idat;
  assign nl_ray_out_rsci_idat = {1'b0 , (ray_out_rsci_idat[164:0])};
  ccs_out_wait_v1 #(.rscid(32'sd62),
  .width(32'sd166)) ray_out_rsci (
      .irdy(ray_out_rsci_irdy),
      .ivld(ray_out_rsci_ivld_hit_sct),
      .idat(nl_ray_out_rsci_idat[165:0]),
      .rdy(ray_out_rsc_rdy),
      .vld(ray_out_rsc_vld),
      .dat(ray_out_rsc_dat)
    );
  WorldHit_hit_ray_out_rsci_ray_out_wait_ctrl WorldHit_hit_ray_out_rsci_ray_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_irdy(ray_out_rsci_irdy),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt),
      .ray_out_rsci_ivld_hit_sct(ray_out_rsci_ivld_hit_sct)
    );
  WorldHit_hit_ray_out_rsci_ray_out_wait_dp WorldHit_hit_ray_out_rsci_ray_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_hit_out_rsci
// ------------------------------------------------------------------


module WorldHit_hit_hit_out_rsci (
  clk, arst_n, hit_out_rsc_dat, hit_out_rsc_vld, hit_out_rsc_rdy, hit_wen, hit_out_rsci_oswt,
      hit_out_rsci_wen_comp, hit_out_rsci_idat
);
  input clk;
  input arst_n;
  output [225:0] hit_out_rsc_dat;
  output hit_out_rsc_vld;
  input hit_out_rsc_rdy;
  input hit_wen;
  input hit_out_rsci_oswt;
  output hit_out_rsci_wen_comp;
  input [225:0] hit_out_rsci_idat;


  // Interconnect Declarations
  wire hit_out_rsci_irdy;
  wire hit_out_rsci_biwt;
  wire hit_out_rsci_bdwt;
  wire hit_out_rsci_bcwt;
  wire hit_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd61),
  .width(32'sd226)) hit_out_rsci (
      .irdy(hit_out_rsci_irdy),
      .ivld(hit_out_rsci_ivld_hit_sct),
      .idat(hit_out_rsci_idat),
      .rdy(hit_out_rsc_rdy),
      .vld(hit_out_rsc_vld),
      .dat(hit_out_rsc_dat)
    );
  WorldHit_hit_hit_out_rsci_hit_out_wait_ctrl WorldHit_hit_hit_out_rsci_hit_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .hit_out_rsci_oswt(hit_out_rsci_oswt),
      .hit_out_rsci_irdy(hit_out_rsci_irdy),
      .hit_out_rsci_biwt(hit_out_rsci_biwt),
      .hit_out_rsci_bdwt(hit_out_rsci_bdwt),
      .hit_out_rsci_bcwt(hit_out_rsci_bcwt),
      .hit_out_rsci_ivld_hit_sct(hit_out_rsci_ivld_hit_sct)
    );
  WorldHit_hit_hit_out_rsci_hit_out_wait_dp WorldHit_hit_hit_out_rsci_hit_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .hit_out_rsci_oswt(hit_out_rsci_oswt),
      .hit_out_rsci_wen_comp(hit_out_rsci_wen_comp),
      .hit_out_rsci_biwt(hit_out_rsci_biwt),
      .hit_out_rsci_bdwt(hit_out_rsci_bdwt),
      .hit_out_rsci_bcwt(hit_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_out_rsci
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_out_rsci (
  clk, arst_n, accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      hit_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  input hit_wen;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input [80:0] accumalated_color_out_rsci_idat;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_irdy;
  wire accumalated_color_out_rsci_biwt;
  wire accumalated_color_out_rsci_bdwt;
  wire accumalated_color_out_rsci_bcwt;
  wire accumalated_color_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd60),
  .width(32'sd81)) accumalated_color_out_rsci (
      .irdy(accumalated_color_out_rsci_irdy),
      .ivld(accumalated_color_out_rsci_ivld_hit_sct),
      .idat(accumalated_color_out_rsci_idat),
      .rdy(accumalated_color_out_rsc_rdy),
      .vld(accumalated_color_out_rsc_vld),
      .dat(accumalated_color_out_rsc_dat)
    );
  WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_irdy(accumalated_color_out_rsci_irdy),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt),
      .accumalated_color_out_rsci_ivld_hit_sct(accumalated_color_out_rsci_ivld_hit_sct)
    );
  WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_dp WorldHit_hit_accumalated_color_out_rsci_accumalated_color_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_out_rsci
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_out_rsci (
  clk, arst_n, attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      hit_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  input hit_wen;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input [80:0] attenuation_chan_out_rsci_idat;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_irdy;
  wire attenuation_chan_out_rsci_biwt;
  wire attenuation_chan_out_rsci_bdwt;
  wire attenuation_chan_out_rsci_bcwt;
  wire attenuation_chan_out_rsci_ivld_hit_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd59),
  .width(32'sd81)) attenuation_chan_out_rsci (
      .irdy(attenuation_chan_out_rsci_irdy),
      .ivld(attenuation_chan_out_rsci_ivld_hit_sct),
      .idat(attenuation_chan_out_rsci_idat),
      .rdy(attenuation_chan_out_rsc_rdy),
      .vld(attenuation_chan_out_rsc_vld),
      .dat(attenuation_chan_out_rsc_dat)
    );
  WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_irdy(attenuation_chan_out_rsci_irdy),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt),
      .attenuation_chan_out_rsci_ivld_hit_sct(attenuation_chan_out_rsci_ivld_hit_sct)
    );
  WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp WorldHit_hit_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outtwo_rsci
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outtwo_rsci (
  clk, arst_n, closest_so_far_outtwo_rsc_dat, closest_so_far_outtwo_rsc_vld, closest_so_far_outtwo_rsc_rdy,
      hit_wen, closest_so_far_outtwo_rsci_oswt, closest_so_far_outtwo_rsci_wen_comp,
      closest_so_far_outtwo_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [46:0] closest_so_far_outtwo_rsc_dat;
  input closest_so_far_outtwo_rsc_vld;
  output closest_so_far_outtwo_rsc_rdy;
  input hit_wen;
  input closest_so_far_outtwo_rsci_oswt;
  output closest_so_far_outtwo_rsci_wen_comp;
  output [46:0] closest_so_far_outtwo_rsci_idat_mxwt;


  // Interconnect Declarations
  wire closest_so_far_outtwo_rsci_biwt;
  wire closest_so_far_outtwo_rsci_bdwt;
  wire closest_so_far_outtwo_rsci_bcwt;
  wire closest_so_far_outtwo_rsci_irdy_hit_sct;
  wire closest_so_far_outtwo_rsci_ivld;
  wire [46:0] closest_so_far_outtwo_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd58),
  .width(32'sd47)) closest_so_far_outtwo_rsci (
      .rdy(closest_so_far_outtwo_rsc_rdy),
      .vld(closest_so_far_outtwo_rsc_vld),
      .dat(closest_so_far_outtwo_rsc_dat),
      .irdy(closest_so_far_outtwo_rsci_irdy_hit_sct),
      .ivld(closest_so_far_outtwo_rsci_ivld),
      .idat(closest_so_far_outtwo_rsci_idat)
    );
  WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_ctrl WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .closest_so_far_outtwo_rsci_oswt(closest_so_far_outtwo_rsci_oswt),
      .closest_so_far_outtwo_rsci_biwt(closest_so_far_outtwo_rsci_biwt),
      .closest_so_far_outtwo_rsci_bdwt(closest_so_far_outtwo_rsci_bdwt),
      .closest_so_far_outtwo_rsci_bcwt(closest_so_far_outtwo_rsci_bcwt),
      .closest_so_far_outtwo_rsci_irdy_hit_sct(closest_so_far_outtwo_rsci_irdy_hit_sct),
      .closest_so_far_outtwo_rsci_ivld(closest_so_far_outtwo_rsci_ivld)
    );
  WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_dp WorldHit_hit_closest_so_far_outtwo_rsci_closest_so_far_outtwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_outtwo_rsci_oswt(closest_so_far_outtwo_rsci_oswt),
      .closest_so_far_outtwo_rsci_wen_comp(closest_so_far_outtwo_rsci_wen_comp),
      .closest_so_far_outtwo_rsci_idat_mxwt(closest_so_far_outtwo_rsci_idat_mxwt),
      .closest_so_far_outtwo_rsci_biwt(closest_so_far_outtwo_rsci_biwt),
      .closest_so_far_outtwo_rsci_bdwt(closest_so_far_outtwo_rsci_bdwt),
      .closest_so_far_outtwo_rsci_bcwt(closest_so_far_outtwo_rsci_bcwt),
      .closest_so_far_outtwo_rsci_idat(closest_so_far_outtwo_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_closest_so_far_outone_rsci
// ------------------------------------------------------------------


module WorldHit_hit_closest_so_far_outone_rsci (
  clk, arst_n, closest_so_far_outone_rsc_dat, closest_so_far_outone_rsc_vld, closest_so_far_outone_rsc_rdy,
      hit_wen, closest_so_far_outone_rsci_oswt, closest_so_far_outone_rsci_wen_comp,
      closest_so_far_outone_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [46:0] closest_so_far_outone_rsc_dat;
  input closest_so_far_outone_rsc_vld;
  output closest_so_far_outone_rsc_rdy;
  input hit_wen;
  input closest_so_far_outone_rsci_oswt;
  output closest_so_far_outone_rsci_wen_comp;
  output [46:0] closest_so_far_outone_rsci_idat_mxwt;


  // Interconnect Declarations
  wire closest_so_far_outone_rsci_biwt;
  wire closest_so_far_outone_rsci_bdwt;
  wire closest_so_far_outone_rsci_bcwt;
  wire closest_so_far_outone_rsci_irdy_hit_sct;
  wire closest_so_far_outone_rsci_ivld;
  wire [46:0] closest_so_far_outone_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd57),
  .width(32'sd47)) closest_so_far_outone_rsci (
      .rdy(closest_so_far_outone_rsc_rdy),
      .vld(closest_so_far_outone_rsc_vld),
      .dat(closest_so_far_outone_rsc_dat),
      .irdy(closest_so_far_outone_rsci_irdy_hit_sct),
      .ivld(closest_so_far_outone_rsci_ivld),
      .idat(closest_so_far_outone_rsci_idat)
    );
  WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_ctrl WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .closest_so_far_outone_rsci_oswt(closest_so_far_outone_rsci_oswt),
      .closest_so_far_outone_rsci_biwt(closest_so_far_outone_rsci_biwt),
      .closest_so_far_outone_rsci_bdwt(closest_so_far_outone_rsci_bdwt),
      .closest_so_far_outone_rsci_bcwt(closest_so_far_outone_rsci_bcwt),
      .closest_so_far_outone_rsci_irdy_hit_sct(closest_so_far_outone_rsci_irdy_hit_sct),
      .closest_so_far_outone_rsci_ivld(closest_so_far_outone_rsci_ivld)
    );
  WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_dp WorldHit_hit_closest_so_far_outone_rsci_closest_so_far_outone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_outone_rsci_oswt(closest_so_far_outone_rsci_oswt),
      .closest_so_far_outone_rsci_wen_comp(closest_so_far_outone_rsci_wen_comp),
      .closest_so_far_outone_rsci_idat_mxwt(closest_so_far_outone_rsci_idat_mxwt),
      .closest_so_far_outone_rsci_biwt(closest_so_far_outone_rsci_biwt),
      .closest_so_far_outone_rsci_bdwt(closest_so_far_outone_rsci_bdwt),
      .closest_so_far_outone_rsci_bcwt(closest_so_far_outone_rsci_bcwt),
      .closest_so_far_outone_rsci_idat(closest_so_far_outone_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outtwo_rsci
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outtwo_rsci (
  clk, arst_n, rec_quad_outtwo_rsc_dat, rec_quad_outtwo_rsc_vld, rec_quad_outtwo_rsc_rdy,
      hit_wen, rec_quad_outtwo_rsci_oswt, rec_quad_outtwo_rsci_wen_comp, rec_quad_outtwo_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [225:0] rec_quad_outtwo_rsc_dat;
  input rec_quad_outtwo_rsc_vld;
  output rec_quad_outtwo_rsc_rdy;
  input hit_wen;
  input rec_quad_outtwo_rsci_oswt;
  output rec_quad_outtwo_rsci_wen_comp;
  output [225:0] rec_quad_outtwo_rsci_idat_mxwt;


  // Interconnect Declarations
  wire rec_quad_outtwo_rsci_biwt;
  wire rec_quad_outtwo_rsci_bdwt;
  wire rec_quad_outtwo_rsci_bcwt;
  wire rec_quad_outtwo_rsci_irdy_hit_sct;
  wire rec_quad_outtwo_rsci_ivld;
  wire [225:0] rec_quad_outtwo_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd56),
  .width(32'sd226)) rec_quad_outtwo_rsci (
      .rdy(rec_quad_outtwo_rsc_rdy),
      .vld(rec_quad_outtwo_rsc_vld),
      .dat(rec_quad_outtwo_rsc_dat),
      .irdy(rec_quad_outtwo_rsci_irdy_hit_sct),
      .ivld(rec_quad_outtwo_rsci_ivld),
      .idat(rec_quad_outtwo_rsci_idat)
    );
  WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_ctrl WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .rec_quad_outtwo_rsci_oswt(rec_quad_outtwo_rsci_oswt),
      .rec_quad_outtwo_rsci_biwt(rec_quad_outtwo_rsci_biwt),
      .rec_quad_outtwo_rsci_bdwt(rec_quad_outtwo_rsci_bdwt),
      .rec_quad_outtwo_rsci_bcwt(rec_quad_outtwo_rsci_bcwt),
      .rec_quad_outtwo_rsci_irdy_hit_sct(rec_quad_outtwo_rsci_irdy_hit_sct),
      .rec_quad_outtwo_rsci_ivld(rec_quad_outtwo_rsci_ivld)
    );
  WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_dp WorldHit_hit_rec_quad_outtwo_rsci_rec_quad_outtwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_outtwo_rsci_oswt(rec_quad_outtwo_rsci_oswt),
      .rec_quad_outtwo_rsci_wen_comp(rec_quad_outtwo_rsci_wen_comp),
      .rec_quad_outtwo_rsci_idat_mxwt(rec_quad_outtwo_rsci_idat_mxwt),
      .rec_quad_outtwo_rsci_biwt(rec_quad_outtwo_rsci_biwt),
      .rec_quad_outtwo_rsci_bdwt(rec_quad_outtwo_rsci_bdwt),
      .rec_quad_outtwo_rsci_bcwt(rec_quad_outtwo_rsci_bcwt),
      .rec_quad_outtwo_rsci_idat(rec_quad_outtwo_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_rec_quad_outone_rsci
// ------------------------------------------------------------------


module WorldHit_hit_rec_quad_outone_rsci (
  clk, arst_n, rec_quad_outone_rsc_dat, rec_quad_outone_rsc_vld, rec_quad_outone_rsc_rdy,
      hit_wen, rec_quad_outone_rsci_oswt, rec_quad_outone_rsci_wen_comp, rec_quad_outone_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [225:0] rec_quad_outone_rsc_dat;
  input rec_quad_outone_rsc_vld;
  output rec_quad_outone_rsc_rdy;
  input hit_wen;
  input rec_quad_outone_rsci_oswt;
  output rec_quad_outone_rsci_wen_comp;
  output [225:0] rec_quad_outone_rsci_idat_mxwt;


  // Interconnect Declarations
  wire rec_quad_outone_rsci_biwt;
  wire rec_quad_outone_rsci_bdwt;
  wire rec_quad_outone_rsci_bcwt;
  wire rec_quad_outone_rsci_irdy_hit_sct;
  wire rec_quad_outone_rsci_ivld;
  wire [225:0] rec_quad_outone_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd55),
  .width(32'sd226)) rec_quad_outone_rsci (
      .rdy(rec_quad_outone_rsc_rdy),
      .vld(rec_quad_outone_rsc_vld),
      .dat(rec_quad_outone_rsc_dat),
      .irdy(rec_quad_outone_rsci_irdy_hit_sct),
      .ivld(rec_quad_outone_rsci_ivld),
      .idat(rec_quad_outone_rsci_idat)
    );
  WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_ctrl WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .rec_quad_outone_rsci_oswt(rec_quad_outone_rsci_oswt),
      .rec_quad_outone_rsci_biwt(rec_quad_outone_rsci_biwt),
      .rec_quad_outone_rsci_bdwt(rec_quad_outone_rsci_bdwt),
      .rec_quad_outone_rsci_bcwt(rec_quad_outone_rsci_bcwt),
      .rec_quad_outone_rsci_irdy_hit_sct(rec_quad_outone_rsci_irdy_hit_sct),
      .rec_quad_outone_rsci_ivld(rec_quad_outone_rsci_ivld)
    );
  WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_dp WorldHit_hit_rec_quad_outone_rsci_rec_quad_outone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_outone_rsci_oswt(rec_quad_outone_rsci_oswt),
      .rec_quad_outone_rsci_wen_comp(rec_quad_outone_rsci_wen_comp),
      .rec_quad_outone_rsci_idat_mxwt(rec_quad_outone_rsci_idat_mxwt),
      .rec_quad_outone_rsci_biwt(rec_quad_outone_rsci_biwt),
      .rec_quad_outone_rsci_bdwt(rec_quad_outone_rsci_bdwt),
      .rec_quad_outone_rsci_bcwt(rec_quad_outone_rsci_bcwt),
      .rec_quad_outone_rsci_idat(rec_quad_outone_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outtwo_rsci
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outtwo_rsci (
  clk, arst_n, quad_hit_anything_outtwo_rsc_dat, quad_hit_anything_outtwo_rsc_vld,
      quad_hit_anything_outtwo_rsc_rdy, hit_wen, quad_hit_anything_outtwo_rsci_oswt,
      quad_hit_anything_outtwo_rsci_wen_comp, quad_hit_anything_outtwo_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input quad_hit_anything_outtwo_rsc_dat;
  input quad_hit_anything_outtwo_rsc_vld;
  output quad_hit_anything_outtwo_rsc_rdy;
  input hit_wen;
  input quad_hit_anything_outtwo_rsci_oswt;
  output quad_hit_anything_outtwo_rsci_wen_comp;
  output quad_hit_anything_outtwo_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quad_hit_anything_outtwo_rsci_biwt;
  wire quad_hit_anything_outtwo_rsci_bdwt;
  wire quad_hit_anything_outtwo_rsci_bcwt;
  wire quad_hit_anything_outtwo_rsci_irdy_hit_sct;
  wire quad_hit_anything_outtwo_rsci_ivld;
  wire quad_hit_anything_outtwo_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd54),
  .width(32'sd1)) quad_hit_anything_outtwo_rsci (
      .rdy(quad_hit_anything_outtwo_rsc_rdy),
      .vld(quad_hit_anything_outtwo_rsc_vld),
      .dat(quad_hit_anything_outtwo_rsc_dat),
      .irdy(quad_hit_anything_outtwo_rsci_irdy_hit_sct),
      .ivld(quad_hit_anything_outtwo_rsci_ivld),
      .idat(quad_hit_anything_outtwo_rsci_idat)
    );
  WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_ctrl WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .quad_hit_anything_outtwo_rsci_oswt(quad_hit_anything_outtwo_rsci_oswt),
      .quad_hit_anything_outtwo_rsci_biwt(quad_hit_anything_outtwo_rsci_biwt),
      .quad_hit_anything_outtwo_rsci_bdwt(quad_hit_anything_outtwo_rsci_bdwt),
      .quad_hit_anything_outtwo_rsci_bcwt(quad_hit_anything_outtwo_rsci_bcwt),
      .quad_hit_anything_outtwo_rsci_irdy_hit_sct(quad_hit_anything_outtwo_rsci_irdy_hit_sct),
      .quad_hit_anything_outtwo_rsci_ivld(quad_hit_anything_outtwo_rsci_ivld)
    );
  WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_dp WorldHit_hit_quad_hit_anything_outtwo_rsci_quad_hit_anything_outtwo_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_outtwo_rsci_oswt(quad_hit_anything_outtwo_rsci_oswt),
      .quad_hit_anything_outtwo_rsci_wen_comp(quad_hit_anything_outtwo_rsci_wen_comp),
      .quad_hit_anything_outtwo_rsci_idat_mxwt(quad_hit_anything_outtwo_rsci_idat_mxwt),
      .quad_hit_anything_outtwo_rsci_biwt(quad_hit_anything_outtwo_rsci_biwt),
      .quad_hit_anything_outtwo_rsci_bdwt(quad_hit_anything_outtwo_rsci_bdwt),
      .quad_hit_anything_outtwo_rsci_bcwt(quad_hit_anything_outtwo_rsci_bcwt),
      .quad_hit_anything_outtwo_rsci_idat(quad_hit_anything_outtwo_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_quad_hit_anything_outone_rsci
// ------------------------------------------------------------------


module WorldHit_hit_quad_hit_anything_outone_rsci (
  clk, arst_n, quad_hit_anything_outone_rsc_dat, quad_hit_anything_outone_rsc_vld,
      quad_hit_anything_outone_rsc_rdy, hit_wen, quad_hit_anything_outone_rsci_oswt,
      quad_hit_anything_outone_rsci_wen_comp, quad_hit_anything_outone_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input quad_hit_anything_outone_rsc_dat;
  input quad_hit_anything_outone_rsc_vld;
  output quad_hit_anything_outone_rsc_rdy;
  input hit_wen;
  input quad_hit_anything_outone_rsci_oswt;
  output quad_hit_anything_outone_rsci_wen_comp;
  output quad_hit_anything_outone_rsci_idat_mxwt;


  // Interconnect Declarations
  wire quad_hit_anything_outone_rsci_biwt;
  wire quad_hit_anything_outone_rsci_bdwt;
  wire quad_hit_anything_outone_rsci_bcwt;
  wire quad_hit_anything_outone_rsci_irdy_hit_sct;
  wire quad_hit_anything_outone_rsci_ivld;
  wire quad_hit_anything_outone_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd53),
  .width(32'sd1)) quad_hit_anything_outone_rsci (
      .rdy(quad_hit_anything_outone_rsc_rdy),
      .vld(quad_hit_anything_outone_rsc_vld),
      .dat(quad_hit_anything_outone_rsc_dat),
      .irdy(quad_hit_anything_outone_rsci_irdy_hit_sct),
      .ivld(quad_hit_anything_outone_rsci_ivld),
      .idat(quad_hit_anything_outone_rsci_idat)
    );
  WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_ctrl WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .quad_hit_anything_outone_rsci_oswt(quad_hit_anything_outone_rsci_oswt),
      .quad_hit_anything_outone_rsci_biwt(quad_hit_anything_outone_rsci_biwt),
      .quad_hit_anything_outone_rsci_bdwt(quad_hit_anything_outone_rsci_bdwt),
      .quad_hit_anything_outone_rsci_bcwt(quad_hit_anything_outone_rsci_bcwt),
      .quad_hit_anything_outone_rsci_irdy_hit_sct(quad_hit_anything_outone_rsci_irdy_hit_sct),
      .quad_hit_anything_outone_rsci_ivld(quad_hit_anything_outone_rsci_ivld)
    );
  WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_dp WorldHit_hit_quad_hit_anything_outone_rsci_quad_hit_anything_outone_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_outone_rsci_oswt(quad_hit_anything_outone_rsci_oswt),
      .quad_hit_anything_outone_rsci_wen_comp(quad_hit_anything_outone_rsci_wen_comp),
      .quad_hit_anything_outone_rsci_idat_mxwt(quad_hit_anything_outone_rsci_idat_mxwt),
      .quad_hit_anything_outone_rsci_biwt(quad_hit_anything_outone_rsci_biwt),
      .quad_hit_anything_outone_rsci_bdwt(quad_hit_anything_outone_rsci_bdwt),
      .quad_hit_anything_outone_rsci_bcwt(quad_hit_anything_outone_rsci_bcwt),
      .quad_hit_anything_outone_rsci_idat(quad_hit_anything_outone_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_accumalated_color_chan_in_rsci
// ------------------------------------------------------------------


module WorldHit_hit_accumalated_color_chan_in_rsci (
  clk, arst_n, accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld,
      accumalated_color_chan_in_rsc_rdy, hit_wen, accumalated_color_chan_in_rsci_oswt,
      accumalated_color_chan_in_rsci_wen_comp, accumalated_color_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input hit_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_biwt;
  wire accumalated_color_chan_in_rsci_bdwt;
  wire accumalated_color_chan_in_rsci_bcwt;
  wire accumalated_color_chan_in_rsci_irdy_hit_sct;
  wire accumalated_color_chan_in_rsci_ivld;
  wire [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd52),
  .width(32'sd81)) accumalated_color_chan_in_rsci (
      .rdy(accumalated_color_chan_in_rsc_rdy),
      .vld(accumalated_color_chan_in_rsc_vld),
      .dat(accumalated_color_chan_in_rsc_dat),
      .irdy(accumalated_color_chan_in_rsci_irdy_hit_sct),
      .ivld(accumalated_color_chan_in_rsci_ivld),
      .idat(accumalated_color_chan_in_rsci_idat)
    );
  WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
      WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_irdy_hit_sct(accumalated_color_chan_in_rsci_irdy_hit_sct),
      .accumalated_color_chan_in_rsci_ivld(accumalated_color_chan_in_rsci_ivld)
    );
  WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp WorldHit_hit_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_idat(accumalated_color_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_attenuation_chan_in_rsci
// ------------------------------------------------------------------


module WorldHit_hit_attenuation_chan_in_rsci (
  clk, arst_n, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      hit_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input hit_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_biwt;
  wire attenuation_chan_in_rsci_bdwt;
  wire attenuation_chan_in_rsci_bcwt;
  wire attenuation_chan_in_rsci_irdy_hit_sct;
  wire attenuation_chan_in_rsci_ivld;
  wire [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd51),
  .width(32'sd81)) attenuation_chan_in_rsci (
      .rdy(attenuation_chan_in_rsc_rdy),
      .vld(attenuation_chan_in_rsc_vld),
      .dat(attenuation_chan_in_rsc_dat),
      .irdy(attenuation_chan_in_rsci_irdy_hit_sct),
      .ivld(attenuation_chan_in_rsci_ivld),
      .idat(attenuation_chan_in_rsci_idat)
    );
  WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_irdy_hit_sct(attenuation_chan_in_rsci_irdy_hit_sct),
      .attenuation_chan_in_rsci_ivld(attenuation_chan_in_rsci_ivld)
    );
  WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp WorldHit_hit_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_idat(attenuation_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_params_in_rsci
// ------------------------------------------------------------------


module WorldHit_hit_params_in_rsci (
  clk, arst_n, params_in_rsc_dat, params_in_rsc_vld, params_in_rsc_rdy, hit_wen,
      params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input hit_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [80:0] params_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire params_in_rsci_biwt;
  wire params_in_rsci_bdwt;
  wire params_in_rsci_bcwt;
  wire params_in_rsci_irdy_hit_sct;
  wire params_in_rsci_ivld;
  wire [92:0] params_in_rsci_idat;
  wire [80:0] params_in_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd50),
  .width(32'sd93)) params_in_rsci (
      .rdy(params_in_rsc_rdy),
      .vld(params_in_rsc_vld),
      .dat(params_in_rsc_dat),
      .irdy(params_in_rsci_irdy_hit_sct),
      .ivld(params_in_rsci_ivld),
      .idat(params_in_rsci_idat)
    );
  WorldHit_hit_params_in_rsci_params_in_wait_ctrl WorldHit_hit_params_in_rsci_params_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_irdy_hit_sct(params_in_rsci_irdy_hit_sct),
      .params_in_rsci_ivld(params_in_rsci_ivld)
    );
  WorldHit_hit_params_in_rsci_params_in_wait_dp WorldHit_hit_params_in_rsci_params_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt_pconst),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_idat(params_in_rsci_idat)
    );
  assign params_in_rsci_idat_mxwt = params_in_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit_ray_in_rsci
// ------------------------------------------------------------------


module WorldHit_hit_ray_in_rsci (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, hit_wen, ray_in_rsci_oswt,
      ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input hit_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [164:0] ray_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_in_rsci_biwt;
  wire ray_in_rsci_bdwt;
  wire ray_in_rsci_bcwt;
  wire ray_in_rsci_irdy_hit_sct;
  wire ray_in_rsci_ivld;
  wire [165:0] ray_in_rsci_idat;
  wire [164:0] ray_in_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd49),
  .width(32'sd166)) ray_in_rsci (
      .rdy(ray_in_rsc_rdy),
      .vld(ray_in_rsc_vld),
      .dat(ray_in_rsc_dat),
      .irdy(ray_in_rsci_irdy_hit_sct),
      .ivld(ray_in_rsci_ivld),
      .idat(ray_in_rsci_idat)
    );
  WorldHit_hit_ray_in_rsci_ray_in_wait_ctrl WorldHit_hit_ray_in_rsci_ray_in_wait_ctrl_inst
      (
      .hit_wen(hit_wen),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_irdy_hit_sct(ray_in_rsci_irdy_hit_sct),
      .ray_in_rsci_ivld(ray_in_rsci_ivld)
    );
  WorldHit_hit_ray_in_rsci_ray_in_wait_dp WorldHit_hit_ray_in_rsci_ray_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt_pconst),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_idat(ray_in_rsci_idat)
    );
  assign ray_in_rsci_idat_mxwt = ray_in_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_out_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_out_rsci (
  clk, arst_n, ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, scatter_wen, ray_out_rsci_oswt,
      ray_out_rsci_wen_comp, ray_out_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  input scatter_wen;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input [165:0] ray_out_rsci_idat;


  // Interconnect Declarations
  wire ray_out_rsci_irdy;
  wire ray_out_rsci_biwt;
  wire ray_out_rsci_bdwt;
  wire ray_out_rsci_bcwt;
  wire ray_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd83),
  .width(32'sd166)) ray_out_rsci (
      .irdy(ray_out_rsci_irdy),
      .ivld(ray_out_rsci_ivld_scatter_sct),
      .idat(ray_out_rsci_idat),
      .rdy(ray_out_rsc_rdy),
      .vld(ray_out_rsc_vld),
      .dat(ray_out_rsc_dat)
    );
  MaterialScatter_scatter_ray_out_rsci_ray_out_wait_ctrl MaterialScatter_scatter_ray_out_rsci_ray_out_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_irdy(ray_out_rsci_irdy),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt),
      .ray_out_rsci_ivld_scatter_sct(ray_out_rsci_ivld_scatter_sct)
    );
  MaterialScatter_scatter_ray_out_rsci_ray_out_wait_dp MaterialScatter_scatter_ray_out_rsci_ray_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_out_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_out_rsci (
  clk, arst_n, accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      scatter_wen, accumalated_color_out_rsci_oswt, accumalated_color_out_rsci_wen_comp,
      accumalated_color_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  input scatter_wen;
  input accumalated_color_out_rsci_oswt;
  output accumalated_color_out_rsci_wen_comp;
  input [80:0] accumalated_color_out_rsci_idat;


  // Interconnect Declarations
  wire accumalated_color_out_rsci_irdy;
  wire accumalated_color_out_rsci_biwt;
  wire accumalated_color_out_rsci_bdwt;
  wire accumalated_color_out_rsci_bcwt;
  wire accumalated_color_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd82),
  .width(32'sd81)) accumalated_color_out_rsci (
      .irdy(accumalated_color_out_rsci_irdy),
      .ivld(accumalated_color_out_rsci_ivld_scatter_sct),
      .idat(accumalated_color_out_rsci_idat),
      .rdy(accumalated_color_out_rsc_rdy),
      .vld(accumalated_color_out_rsc_vld),
      .dat(accumalated_color_out_rsc_dat)
    );
  MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl
      MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_irdy(accumalated_color_out_rsci_irdy),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt),
      .accumalated_color_out_rsci_ivld_scatter_sct(accumalated_color_out_rsci_ivld_scatter_sct)
    );
  MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_dp
      MaterialScatter_scatter_accumalated_color_out_rsci_accumalated_color_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsci_oswt(accumalated_color_out_rsci_oswt),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_biwt(accumalated_color_out_rsci_biwt),
      .accumalated_color_out_rsci_bdwt(accumalated_color_out_rsci_bdwt),
      .accumalated_color_out_rsci_bcwt(accumalated_color_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_out_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_out_rsci (
  clk, arst_n, attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      scatter_wen, attenuation_chan_out_rsci_oswt, attenuation_chan_out_rsci_wen_comp,
      attenuation_chan_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  input scatter_wen;
  input attenuation_chan_out_rsci_oswt;
  output attenuation_chan_out_rsci_wen_comp;
  input [80:0] attenuation_chan_out_rsci_idat;


  // Interconnect Declarations
  wire attenuation_chan_out_rsci_irdy;
  wire attenuation_chan_out_rsci_biwt;
  wire attenuation_chan_out_rsci_bdwt;
  wire attenuation_chan_out_rsci_bcwt;
  wire attenuation_chan_out_rsci_ivld_scatter_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd81),
  .width(32'sd81)) attenuation_chan_out_rsci (
      .irdy(attenuation_chan_out_rsci_irdy),
      .ivld(attenuation_chan_out_rsci_ivld_scatter_sct),
      .idat(attenuation_chan_out_rsci_idat),
      .rdy(attenuation_chan_out_rsc_rdy),
      .vld(attenuation_chan_out_rsc_vld),
      .dat(attenuation_chan_out_rsc_dat)
    );
  MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl
      MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_irdy(attenuation_chan_out_rsci_irdy),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt),
      .attenuation_chan_out_rsci_ivld_scatter_sct(attenuation_chan_out_rsci_ivld_scatter_sct)
    );
  MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp
      MaterialScatter_scatter_attenuation_chan_out_rsci_attenuation_chan_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsci_oswt(attenuation_chan_out_rsci_oswt),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_biwt(attenuation_chan_out_rsci_biwt),
      .attenuation_chan_out_rsci_bdwt(attenuation_chan_out_rsci_bdwt),
      .attenuation_chan_out_rsci_bcwt(attenuation_chan_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_isHit_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_isHit_rsci (
  clk, arst_n, isHit_rsc_dat, isHit_rsc_vld, isHit_rsc_rdy, scatter_wen, isHit_rsci_oswt,
      isHit_rsci_wen_comp, isHit_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input isHit_rsc_dat;
  input isHit_rsc_vld;
  output isHit_rsc_rdy;
  input scatter_wen;
  input isHit_rsci_oswt;
  output isHit_rsci_wen_comp;
  output isHit_rsci_idat_mxwt;


  // Interconnect Declarations
  wire isHit_rsci_biwt;
  wire isHit_rsci_bdwt;
  wire isHit_rsci_bcwt;
  wire isHit_rsci_irdy_scatter_sct;
  wire isHit_rsci_ivld;
  wire isHit_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd80),
  .width(32'sd1)) isHit_rsci (
      .rdy(isHit_rsc_rdy),
      .vld(isHit_rsc_vld),
      .dat(isHit_rsc_dat),
      .irdy(isHit_rsci_irdy_scatter_sct),
      .ivld(isHit_rsci_ivld),
      .idat(isHit_rsci_idat)
    );
  MaterialScatter_scatter_isHit_rsci_isHit_wait_ctrl MaterialScatter_scatter_isHit_rsci_isHit_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .isHit_rsci_oswt(isHit_rsci_oswt),
      .isHit_rsci_biwt(isHit_rsci_biwt),
      .isHit_rsci_bdwt(isHit_rsci_bdwt),
      .isHit_rsci_bcwt(isHit_rsci_bcwt),
      .isHit_rsci_irdy_scatter_sct(isHit_rsci_irdy_scatter_sct),
      .isHit_rsci_ivld(isHit_rsci_ivld)
    );
  MaterialScatter_scatter_isHit_rsci_isHit_wait_dp MaterialScatter_scatter_isHit_rsci_isHit_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .isHit_rsci_oswt(isHit_rsci_oswt),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp),
      .isHit_rsci_idat_mxwt(isHit_rsci_idat_mxwt),
      .isHit_rsci_biwt(isHit_rsci_biwt),
      .isHit_rsci_bdwt(isHit_rsci_bdwt),
      .isHit_rsci_bcwt(isHit_rsci_bcwt),
      .isHit_rsci_idat(isHit_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_accumalated_color_chan_in_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_accumalated_color_chan_in_rsci (
  clk, arst_n, accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld,
      accumalated_color_chan_in_rsc_rdy, scatter_wen, accumalated_color_chan_in_rsci_oswt,
      accumalated_color_chan_in_rsci_wen_comp, accumalated_color_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input scatter_wen;
  input accumalated_color_chan_in_rsci_oswt;
  output accumalated_color_chan_in_rsci_wen_comp;
  output [80:0] accumalated_color_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire accumalated_color_chan_in_rsci_biwt;
  wire accumalated_color_chan_in_rsci_bdwt;
  wire accumalated_color_chan_in_rsci_bcwt;
  wire accumalated_color_chan_in_rsci_irdy_scatter_sct;
  wire accumalated_color_chan_in_rsci_ivld;
  wire [80:0] accumalated_color_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd79),
  .width(32'sd81)) accumalated_color_chan_in_rsci (
      .rdy(accumalated_color_chan_in_rsc_rdy),
      .vld(accumalated_color_chan_in_rsc_vld),
      .dat(accumalated_color_chan_in_rsc_dat),
      .irdy(accumalated_color_chan_in_rsci_irdy_scatter_sct),
      .ivld(accumalated_color_chan_in_rsci_ivld),
      .idat(accumalated_color_chan_in_rsci_idat)
    );
  MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl
      MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_irdy_scatter_sct(accumalated_color_chan_in_rsci_irdy_scatter_sct),
      .accumalated_color_chan_in_rsci_ivld(accumalated_color_chan_in_rsci_ivld)
    );
  MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp
      MaterialScatter_scatter_accumalated_color_chan_in_rsci_accumalated_color_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsci_oswt(accumalated_color_chan_in_rsci_oswt),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt),
      .accumalated_color_chan_in_rsci_biwt(accumalated_color_chan_in_rsci_biwt),
      .accumalated_color_chan_in_rsci_bdwt(accumalated_color_chan_in_rsci_bdwt),
      .accumalated_color_chan_in_rsci_bcwt(accumalated_color_chan_in_rsci_bcwt),
      .accumalated_color_chan_in_rsci_idat(accumalated_color_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_attenuation_chan_in_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_attenuation_chan_in_rsci (
  clk, arst_n, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      scatter_wen, attenuation_chan_in_rsci_oswt, attenuation_chan_in_rsci_wen_comp,
      attenuation_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input scatter_wen;
  input attenuation_chan_in_rsci_oswt;
  output attenuation_chan_in_rsci_wen_comp;
  output [80:0] attenuation_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire attenuation_chan_in_rsci_biwt;
  wire attenuation_chan_in_rsci_bdwt;
  wire attenuation_chan_in_rsci_bcwt;
  wire attenuation_chan_in_rsci_irdy_scatter_sct;
  wire attenuation_chan_in_rsci_ivld;
  wire [80:0] attenuation_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd78),
  .width(32'sd81)) attenuation_chan_in_rsci (
      .rdy(attenuation_chan_in_rsc_rdy),
      .vld(attenuation_chan_in_rsc_vld),
      .dat(attenuation_chan_in_rsc_dat),
      .irdy(attenuation_chan_in_rsci_irdy_scatter_sct),
      .ivld(attenuation_chan_in_rsci_ivld),
      .idat(attenuation_chan_in_rsci_idat)
    );
  MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl
      MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_irdy_scatter_sct(attenuation_chan_in_rsci_irdy_scatter_sct),
      .attenuation_chan_in_rsci_ivld(attenuation_chan_in_rsci_ivld)
    );
  MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp MaterialScatter_scatter_attenuation_chan_in_rsci_attenuation_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsci_oswt(attenuation_chan_in_rsci_oswt),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt),
      .attenuation_chan_in_rsci_biwt(attenuation_chan_in_rsci_biwt),
      .attenuation_chan_in_rsci_bdwt(attenuation_chan_in_rsci_bdwt),
      .attenuation_chan_in_rsci_bcwt(attenuation_chan_in_rsci_bcwt),
      .attenuation_chan_in_rsci_idat(attenuation_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_hit_in_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_hit_in_rsci (
  clk, arst_n, hit_in_rsc_dat, hit_in_rsc_vld, hit_in_rsc_rdy, scatter_wen, hit_in_rsci_oswt,
      hit_in_rsci_wen_comp, hit_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [225:0] hit_in_rsc_dat;
  input hit_in_rsc_vld;
  output hit_in_rsc_rdy;
  input scatter_wen;
  input hit_in_rsci_oswt;
  output hit_in_rsci_wen_comp;
  output [225:0] hit_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire hit_in_rsci_biwt;
  wire hit_in_rsci_bdwt;
  wire hit_in_rsci_bcwt;
  wire hit_in_rsci_irdy_scatter_sct;
  wire hit_in_rsci_ivld;
  wire [225:0] hit_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd77),
  .width(32'sd226)) hit_in_rsci (
      .rdy(hit_in_rsc_rdy),
      .vld(hit_in_rsc_vld),
      .dat(hit_in_rsc_dat),
      .irdy(hit_in_rsci_irdy_scatter_sct),
      .ivld(hit_in_rsci_ivld),
      .idat(hit_in_rsci_idat)
    );
  MaterialScatter_scatter_hit_in_rsci_hit_in_wait_ctrl MaterialScatter_scatter_hit_in_rsci_hit_in_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .hit_in_rsci_oswt(hit_in_rsci_oswt),
      .hit_in_rsci_biwt(hit_in_rsci_biwt),
      .hit_in_rsci_bdwt(hit_in_rsci_bdwt),
      .hit_in_rsci_bcwt(hit_in_rsci_bcwt),
      .hit_in_rsci_irdy_scatter_sct(hit_in_rsci_irdy_scatter_sct),
      .hit_in_rsci_ivld(hit_in_rsci_ivld)
    );
  MaterialScatter_scatter_hit_in_rsci_hit_in_wait_dp MaterialScatter_scatter_hit_in_rsci_hit_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .hit_in_rsci_oswt(hit_in_rsci_oswt),
      .hit_in_rsci_wen_comp(hit_in_rsci_wen_comp),
      .hit_in_rsci_idat_mxwt(hit_in_rsci_idat_mxwt),
      .hit_in_rsci_biwt(hit_in_rsci_biwt),
      .hit_in_rsci_bdwt(hit_in_rsci_bdwt),
      .hit_in_rsci_bcwt(hit_in_rsci_bcwt),
      .hit_in_rsci_idat(hit_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter_ray_in_rsci
// ------------------------------------------------------------------


module MaterialScatter_scatter_ray_in_rsci (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, scatter_wen, ray_in_rsci_oswt,
      ray_in_rsci_wen_comp, ray_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input scatter_wen;
  input ray_in_rsci_oswt;
  output ray_in_rsci_wen_comp;
  output [165:0] ray_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_in_rsci_biwt;
  wire ray_in_rsci_bdwt;
  wire ray_in_rsci_bcwt;
  wire ray_in_rsci_irdy_scatter_sct;
  wire ray_in_rsci_ivld;
  wire [165:0] ray_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd76),
  .width(32'sd166)) ray_in_rsci (
      .rdy(ray_in_rsc_rdy),
      .vld(ray_in_rsc_vld),
      .dat(ray_in_rsc_dat),
      .irdy(ray_in_rsci_irdy_scatter_sct),
      .ivld(ray_in_rsci_ivld),
      .idat(ray_in_rsci_idat)
    );
  MaterialScatter_scatter_ray_in_rsci_ray_in_wait_ctrl MaterialScatter_scatter_ray_in_rsci_ray_in_wait_ctrl_inst
      (
      .scatter_wen(scatter_wen),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_irdy_scatter_sct(ray_in_rsci_irdy_scatter_sct),
      .ray_in_rsci_ivld(ray_in_rsci_ivld)
    );
  MaterialScatter_scatter_ray_in_rsci_ray_in_wait_dp MaterialScatter_scatter_ray_in_rsci_ray_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsci_oswt(ray_in_rsci_oswt),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt),
      .ray_in_rsci_biwt(ray_in_rsci_biwt),
      .ray_in_rsci_bdwt(ray_in_rsci_bdwt),
      .ray_in_rsci_bcwt(ray_in_rsci_bcwt),
      .ray_in_rsci_idat(ray_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_output_pxl_serial_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_output_pxl_serial_rsci (
  clk, arst_n, output_pxl_serial_rsc_dat, output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy,
      run_wen, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_wen_comp, output_pxl_serial_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;
  input run_wen;
  input output_pxl_serial_rsci_oswt;
  output output_pxl_serial_rsci_wen_comp;
  input [80:0] output_pxl_serial_rsci_idat;


  // Interconnect Declarations
  wire output_pxl_serial_rsci_irdy;
  wire output_pxl_serial_rsci_biwt;
  wire output_pxl_serial_rsci_bdwt;
  wire output_pxl_serial_rsci_bcwt;
  wire output_pxl_serial_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd124),
  .width(32'sd81)) output_pxl_serial_rsci (
      .irdy(output_pxl_serial_rsci_irdy),
      .ivld(output_pxl_serial_rsci_ivld_run_sct),
      .idat(output_pxl_serial_rsci_idat),
      .rdy(output_pxl_serial_rsc_rdy),
      .vld(output_pxl_serial_rsc_vld),
      .dat(output_pxl_serial_rsc_dat)
    );
  ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl
      ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .output_pxl_serial_rsci_oswt(output_pxl_serial_rsci_oswt),
      .output_pxl_serial_rsci_irdy(output_pxl_serial_rsci_irdy),
      .output_pxl_serial_rsci_biwt(output_pxl_serial_rsci_biwt),
      .output_pxl_serial_rsci_bdwt(output_pxl_serial_rsci_bdwt),
      .output_pxl_serial_rsci_bcwt(output_pxl_serial_rsci_bcwt),
      .output_pxl_serial_rsci_ivld_run_sct(output_pxl_serial_rsci_ivld_run_sct)
    );
  ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp ShaderFeedbackController_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_pxl_serial_rsci_oswt(output_pxl_serial_rsci_oswt),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp),
      .output_pxl_serial_rsci_biwt(output_pxl_serial_rsci_biwt),
      .output_pxl_serial_rsci_bdwt(output_pxl_serial_rsci_bdwt),
      .output_pxl_serial_rsci_bcwt(output_pxl_serial_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_out_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_out_rsci (
  clk, arst_n, atten_chan_out_rsc_dat, atten_chan_out_rsc_vld, atten_chan_out_rsc_rdy,
      run_wen, atten_chan_out_rsci_oswt, atten_chan_out_rsci_wen_comp, atten_chan_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] atten_chan_out_rsc_dat;
  output atten_chan_out_rsc_vld;
  input atten_chan_out_rsc_rdy;
  input run_wen;
  input atten_chan_out_rsci_oswt;
  output atten_chan_out_rsci_wen_comp;
  input [80:0] atten_chan_out_rsci_idat;


  // Interconnect Declarations
  wire atten_chan_out_rsci_irdy;
  wire atten_chan_out_rsci_biwt;
  wire atten_chan_out_rsci_bdwt;
  wire atten_chan_out_rsci_bcwt;
  wire atten_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd123),
  .width(32'sd81)) atten_chan_out_rsci (
      .irdy(atten_chan_out_rsci_irdy),
      .ivld(atten_chan_out_rsci_ivld_run_sct),
      .idat(atten_chan_out_rsci_idat),
      .rdy(atten_chan_out_rsc_rdy),
      .vld(atten_chan_out_rsc_vld),
      .dat(atten_chan_out_rsc_dat)
    );
  ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_ctrl ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .atten_chan_out_rsci_oswt(atten_chan_out_rsci_oswt),
      .atten_chan_out_rsci_irdy(atten_chan_out_rsci_irdy),
      .atten_chan_out_rsci_biwt(atten_chan_out_rsci_biwt),
      .atten_chan_out_rsci_bdwt(atten_chan_out_rsci_bdwt),
      .atten_chan_out_rsci_bcwt(atten_chan_out_rsci_bcwt),
      .atten_chan_out_rsci_ivld_run_sct(atten_chan_out_rsci_ivld_run_sct)
    );
  ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_dp ShaderFeedbackController_run_atten_chan_out_rsci_atten_chan_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .atten_chan_out_rsci_oswt(atten_chan_out_rsci_oswt),
      .atten_chan_out_rsci_wen_comp(atten_chan_out_rsci_wen_comp),
      .atten_chan_out_rsci_biwt(atten_chan_out_rsci_biwt),
      .atten_chan_out_rsci_bdwt(atten_chan_out_rsci_bdwt),
      .atten_chan_out_rsci_bcwt(atten_chan_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_out_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_out_rsci (
  clk, arst_n, color_chan_out_rsc_dat, color_chan_out_rsc_vld, color_chan_out_rsc_rdy,
      run_wen, color_chan_out_rsci_oswt, color_chan_out_rsci_wen_comp, color_chan_out_rsci_idat
);
  input clk;
  input arst_n;
  output [80:0] color_chan_out_rsc_dat;
  output color_chan_out_rsc_vld;
  input color_chan_out_rsc_rdy;
  input run_wen;
  input color_chan_out_rsci_oswt;
  output color_chan_out_rsci_wen_comp;
  input [80:0] color_chan_out_rsci_idat;


  // Interconnect Declarations
  wire color_chan_out_rsci_irdy;
  wire color_chan_out_rsci_biwt;
  wire color_chan_out_rsci_bdwt;
  wire color_chan_out_rsci_bcwt;
  wire color_chan_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd122),
  .width(32'sd81)) color_chan_out_rsci (
      .irdy(color_chan_out_rsci_irdy),
      .ivld(color_chan_out_rsci_ivld_run_sct),
      .idat(color_chan_out_rsci_idat),
      .rdy(color_chan_out_rsc_rdy),
      .vld(color_chan_out_rsc_vld),
      .dat(color_chan_out_rsc_dat)
    );
  ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_ctrl ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .color_chan_out_rsci_oswt(color_chan_out_rsci_oswt),
      .color_chan_out_rsci_irdy(color_chan_out_rsci_irdy),
      .color_chan_out_rsci_biwt(color_chan_out_rsci_biwt),
      .color_chan_out_rsci_bdwt(color_chan_out_rsci_bdwt),
      .color_chan_out_rsci_bcwt(color_chan_out_rsci_bcwt),
      .color_chan_out_rsci_ivld_run_sct(color_chan_out_rsci_ivld_run_sct)
    );
  ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_dp ShaderFeedbackController_run_color_chan_out_rsci_color_chan_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .color_chan_out_rsci_oswt(color_chan_out_rsci_oswt),
      .color_chan_out_rsci_wen_comp(color_chan_out_rsci_wen_comp),
      .color_chan_out_rsci_biwt(color_chan_out_rsci_biwt),
      .color_chan_out_rsci_bdwt(color_chan_out_rsci_bdwt),
      .color_chan_out_rsci_bcwt(color_chan_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_out_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_out_rsci (
  clk, arst_n, params_out_rsc_dat, params_out_rsc_vld, params_out_rsc_rdy, run_wen,
      params_out_rsci_oswt, params_out_rsci_wen_comp, params_out_rsci_idat
);
  input clk;
  input arst_n;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;
  input run_wen;
  input params_out_rsci_oswt;
  output params_out_rsci_wen_comp;
  input [92:0] params_out_rsci_idat;


  // Interconnect Declarations
  wire params_out_rsci_irdy;
  wire params_out_rsci_biwt;
  wire params_out_rsci_bdwt;
  wire params_out_rsci_bcwt;
  wire params_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd121),
  .width(32'sd93)) params_out_rsci (
      .irdy(params_out_rsci_irdy),
      .ivld(params_out_rsci_ivld_run_sct),
      .idat(params_out_rsci_idat),
      .rdy(params_out_rsc_rdy),
      .vld(params_out_rsc_vld),
      .dat(params_out_rsc_dat)
    );
  ShaderFeedbackController_run_params_out_rsci_params_out_wait_ctrl ShaderFeedbackController_run_params_out_rsci_params_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .params_out_rsci_oswt(params_out_rsci_oswt),
      .params_out_rsci_irdy(params_out_rsci_irdy),
      .params_out_rsci_biwt(params_out_rsci_biwt),
      .params_out_rsci_bdwt(params_out_rsci_bdwt),
      .params_out_rsci_bcwt(params_out_rsci_bcwt),
      .params_out_rsci_ivld_run_sct(params_out_rsci_ivld_run_sct)
    );
  ShaderFeedbackController_run_params_out_rsci_params_out_wait_dp ShaderFeedbackController_run_params_out_rsci_params_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_out_rsci_oswt(params_out_rsci_oswt),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp),
      .params_out_rsci_biwt(params_out_rsci_biwt),
      .params_out_rsci_bdwt(params_out_rsci_bdwt),
      .params_out_rsci_bcwt(params_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_out_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_out_rsci (
  clk, arst_n, ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, run_wen, ray_out_rsci_oswt,
      ray_out_rsci_wen_comp, ray_out_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  input run_wen;
  input ray_out_rsci_oswt;
  output ray_out_rsci_wen_comp;
  input [165:0] ray_out_rsci_idat;


  // Interconnect Declarations
  wire ray_out_rsci_irdy;
  wire ray_out_rsci_biwt;
  wire ray_out_rsci_bdwt;
  wire ray_out_rsci_bcwt;
  wire ray_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd120),
  .width(32'sd166)) ray_out_rsci (
      .irdy(ray_out_rsci_irdy),
      .ivld(ray_out_rsci_ivld_run_sct),
      .idat(ray_out_rsci_idat),
      .rdy(ray_out_rsc_rdy),
      .vld(ray_out_rsc_vld),
      .dat(ray_out_rsc_dat)
    );
  ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_ctrl ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_irdy(ray_out_rsci_irdy),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt),
      .ray_out_rsci_ivld_run_sct(ray_out_rsci_ivld_run_sct)
    );
  ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_dp ShaderFeedbackController_run_ray_out_rsci_ray_out_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsci_oswt(ray_out_rsci_oswt),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_biwt(ray_out_rsci_biwt),
      .ray_out_rsci_bdwt(ray_out_rsci_bdwt),
      .ray_out_rsci_bcwt(ray_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_atten_chan_in_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_atten_chan_in_rsci (
  clk, arst_n, atten_chan_in_rsc_dat, atten_chan_in_rsc_vld, atten_chan_in_rsc_rdy,
      run_wen, atten_chan_in_rsci_oswt, atten_chan_in_rsci_wen_comp, atten_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] atten_chan_in_rsc_dat;
  input atten_chan_in_rsc_vld;
  output atten_chan_in_rsc_rdy;
  input run_wen;
  input atten_chan_in_rsci_oswt;
  output atten_chan_in_rsci_wen_comp;
  output [80:0] atten_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire atten_chan_in_rsci_biwt;
  wire atten_chan_in_rsci_bdwt;
  wire atten_chan_in_rsci_bcwt;
  wire atten_chan_in_rsci_irdy_run_sct;
  wire atten_chan_in_rsci_ivld;
  wire [80:0] atten_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd119),
  .width(32'sd81)) atten_chan_in_rsci (
      .rdy(atten_chan_in_rsc_rdy),
      .vld(atten_chan_in_rsc_vld),
      .dat(atten_chan_in_rsc_dat),
      .irdy(atten_chan_in_rsci_irdy_run_sct),
      .ivld(atten_chan_in_rsci_ivld),
      .idat(atten_chan_in_rsci_idat)
    );
  ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_ctrl ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .atten_chan_in_rsci_oswt(atten_chan_in_rsci_oswt),
      .atten_chan_in_rsci_biwt(atten_chan_in_rsci_biwt),
      .atten_chan_in_rsci_bdwt(atten_chan_in_rsci_bdwt),
      .atten_chan_in_rsci_bcwt(atten_chan_in_rsci_bcwt),
      .atten_chan_in_rsci_irdy_run_sct(atten_chan_in_rsci_irdy_run_sct),
      .atten_chan_in_rsci_ivld(atten_chan_in_rsci_ivld)
    );
  ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_dp ShaderFeedbackController_run_atten_chan_in_rsci_atten_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .atten_chan_in_rsci_oswt(atten_chan_in_rsci_oswt),
      .atten_chan_in_rsci_wen_comp(atten_chan_in_rsci_wen_comp),
      .atten_chan_in_rsci_idat_mxwt(atten_chan_in_rsci_idat_mxwt),
      .atten_chan_in_rsci_biwt(atten_chan_in_rsci_biwt),
      .atten_chan_in_rsci_bdwt(atten_chan_in_rsci_bdwt),
      .atten_chan_in_rsci_bcwt(atten_chan_in_rsci_bcwt),
      .atten_chan_in_rsci_idat(atten_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_color_chan_in_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_color_chan_in_rsci (
  clk, arst_n, color_chan_in_rsc_dat, color_chan_in_rsc_vld, color_chan_in_rsc_rdy,
      run_wen, color_chan_in_rsci_oswt, color_chan_in_rsci_wen_comp, color_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] color_chan_in_rsc_dat;
  input color_chan_in_rsc_vld;
  output color_chan_in_rsc_rdy;
  input run_wen;
  input color_chan_in_rsci_oswt;
  output color_chan_in_rsci_wen_comp;
  output [80:0] color_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire color_chan_in_rsci_biwt;
  wire color_chan_in_rsci_bdwt;
  wire color_chan_in_rsci_bcwt;
  wire color_chan_in_rsci_irdy_run_sct;
  wire color_chan_in_rsci_ivld;
  wire [80:0] color_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd118),
  .width(32'sd81)) color_chan_in_rsci (
      .rdy(color_chan_in_rsc_rdy),
      .vld(color_chan_in_rsc_vld),
      .dat(color_chan_in_rsc_dat),
      .irdy(color_chan_in_rsci_irdy_run_sct),
      .ivld(color_chan_in_rsci_ivld),
      .idat(color_chan_in_rsci_idat)
    );
  ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_ctrl ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .color_chan_in_rsci_oswt(color_chan_in_rsci_oswt),
      .color_chan_in_rsci_biwt(color_chan_in_rsci_biwt),
      .color_chan_in_rsci_bdwt(color_chan_in_rsci_bdwt),
      .color_chan_in_rsci_bcwt(color_chan_in_rsci_bcwt),
      .color_chan_in_rsci_irdy_run_sct(color_chan_in_rsci_irdy_run_sct),
      .color_chan_in_rsci_ivld(color_chan_in_rsci_ivld)
    );
  ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_dp ShaderFeedbackController_run_color_chan_in_rsci_color_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .color_chan_in_rsci_oswt(color_chan_in_rsci_oswt),
      .color_chan_in_rsci_wen_comp(color_chan_in_rsci_wen_comp),
      .color_chan_in_rsci_idat_mxwt(color_chan_in_rsci_idat_mxwt),
      .color_chan_in_rsci_biwt(color_chan_in_rsci_biwt),
      .color_chan_in_rsci_bdwt(color_chan_in_rsci_bdwt),
      .color_chan_in_rsci_bcwt(color_chan_in_rsci_bcwt),
      .color_chan_in_rsci_idat(color_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_params_in_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_params_in_rsci (
  clk, arst_n, params_in_rsc_dat, params_in_rsc_vld, params_in_rsc_rdy, run_wen,
      params_in_rsci_oswt, params_in_rsci_wen_comp, params_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input run_wen;
  input params_in_rsci_oswt;
  output params_in_rsci_wen_comp;
  output [92:0] params_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire params_in_rsci_biwt;
  wire params_in_rsci_bdwt;
  wire params_in_rsci_bcwt;
  wire params_in_rsci_irdy_run_sct;
  wire params_in_rsci_ivld;
  wire [92:0] params_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd117),
  .width(32'sd93)) params_in_rsci (
      .rdy(params_in_rsc_rdy),
      .vld(params_in_rsc_vld),
      .dat(params_in_rsc_dat),
      .irdy(params_in_rsci_irdy_run_sct),
      .ivld(params_in_rsci_ivld),
      .idat(params_in_rsci_idat)
    );
  ShaderFeedbackController_run_params_in_rsci_params_in_wait_ctrl ShaderFeedbackController_run_params_in_rsci_params_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_irdy_run_sct(params_in_rsci_irdy_run_sct),
      .params_in_rsci_ivld(params_in_rsci_ivld)
    );
  ShaderFeedbackController_run_params_in_rsci_params_in_wait_dp ShaderFeedbackController_run_params_in_rsci_params_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsci_oswt(params_in_rsci_oswt),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt),
      .params_in_rsci_biwt(params_in_rsci_biwt),
      .params_in_rsci_bdwt(params_in_rsci_bdwt),
      .params_in_rsci_bcwt(params_in_rsci_bcwt),
      .params_in_rsci_idat(params_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_scattered_chan_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_scattered_chan_rsci (
  clk, arst_n, ray_scattered_chan_rsc_dat, ray_scattered_chan_rsc_vld, ray_scattered_chan_rsc_rdy,
      run_wen, ray_scattered_chan_rsci_oswt, ray_scattered_chan_rsci_wen_comp, ray_scattered_chan_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_scattered_chan_rsc_dat;
  input ray_scattered_chan_rsc_vld;
  output ray_scattered_chan_rsc_rdy;
  input run_wen;
  input ray_scattered_chan_rsci_oswt;
  output ray_scattered_chan_rsci_wen_comp;
  output [165:0] ray_scattered_chan_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_scattered_chan_rsci_biwt;
  wire ray_scattered_chan_rsci_bdwt;
  wire ray_scattered_chan_rsci_bcwt;
  wire ray_scattered_chan_rsci_irdy_run_sct;
  wire ray_scattered_chan_rsci_ivld;
  wire [165:0] ray_scattered_chan_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd116),
  .width(32'sd166)) ray_scattered_chan_rsci (
      .rdy(ray_scattered_chan_rsc_rdy),
      .vld(ray_scattered_chan_rsc_vld),
      .dat(ray_scattered_chan_rsc_dat),
      .irdy(ray_scattered_chan_rsci_irdy_run_sct),
      .ivld(ray_scattered_chan_rsci_ivld),
      .idat(ray_scattered_chan_rsci_idat)
    );
  ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_ctrl
      ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_scattered_chan_rsci_oswt(ray_scattered_chan_rsci_oswt),
      .ray_scattered_chan_rsci_biwt(ray_scattered_chan_rsci_biwt),
      .ray_scattered_chan_rsci_bdwt(ray_scattered_chan_rsci_bdwt),
      .ray_scattered_chan_rsci_bcwt(ray_scattered_chan_rsci_bcwt),
      .ray_scattered_chan_rsci_irdy_run_sct(ray_scattered_chan_rsci_irdy_run_sct),
      .ray_scattered_chan_rsci_ivld(ray_scattered_chan_rsci_ivld)
    );
  ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_dp
      ShaderFeedbackController_run_ray_scattered_chan_rsci_ray_scattered_chan_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_scattered_chan_rsci_oswt(ray_scattered_chan_rsci_oswt),
      .ray_scattered_chan_rsci_wen_comp(ray_scattered_chan_rsci_wen_comp),
      .ray_scattered_chan_rsci_idat_mxwt(ray_scattered_chan_rsci_idat_mxwt),
      .ray_scattered_chan_rsci_biwt(ray_scattered_chan_rsci_biwt),
      .ray_scattered_chan_rsci_bdwt(ray_scattered_chan_rsci_bdwt),
      .ray_scattered_chan_rsci_bcwt(ray_scattered_chan_rsci_bcwt),
      .ray_scattered_chan_rsci_idat(ray_scattered_chan_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run_ray_chan_in_rsci
// ------------------------------------------------------------------


module ShaderFeedbackController_run_ray_chan_in_rsci (
  clk, arst_n, ray_chan_in_rsc_dat, ray_chan_in_rsc_vld, ray_chan_in_rsc_rdy, run_wen,
      ray_chan_in_rsci_oswt, ray_chan_in_rsci_wen_comp, ray_chan_in_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] ray_chan_in_rsc_dat;
  input ray_chan_in_rsc_vld;
  output ray_chan_in_rsc_rdy;
  input run_wen;
  input ray_chan_in_rsci_oswt;
  output ray_chan_in_rsci_wen_comp;
  output [165:0] ray_chan_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ray_chan_in_rsci_biwt;
  wire ray_chan_in_rsci_bdwt;
  wire ray_chan_in_rsci_bcwt;
  wire ray_chan_in_rsci_irdy_run_sct;
  wire ray_chan_in_rsci_ivld;
  wire [165:0] ray_chan_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd115),
  .width(32'sd166)) ray_chan_in_rsci (
      .rdy(ray_chan_in_rsc_rdy),
      .vld(ray_chan_in_rsc_vld),
      .dat(ray_chan_in_rsc_dat),
      .irdy(ray_chan_in_rsci_irdy_run_sct),
      .ivld(ray_chan_in_rsci_ivld),
      .idat(ray_chan_in_rsci_idat)
    );
  ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_ctrl ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ray_chan_in_rsci_oswt(ray_chan_in_rsci_oswt),
      .ray_chan_in_rsci_biwt(ray_chan_in_rsci_biwt),
      .ray_chan_in_rsci_bdwt(ray_chan_in_rsci_bdwt),
      .ray_chan_in_rsci_bcwt(ray_chan_in_rsci_bcwt),
      .ray_chan_in_rsci_irdy_run_sct(ray_chan_in_rsci_irdy_run_sct),
      .ray_chan_in_rsci_ivld(ray_chan_in_rsci_ivld)
    );
  ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_dp ShaderFeedbackController_run_ray_chan_in_rsci_ray_chan_in_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_chan_in_rsci_oswt(ray_chan_in_rsci_oswt),
      .ray_chan_in_rsci_wen_comp(ray_chan_in_rsci_wen_comp),
      .ray_chan_in_rsci_idat_mxwt(ray_chan_in_rsci_idat_mxwt),
      .ray_chan_in_rsci_biwt(ray_chan_in_rsci_biwt),
      .ray_chan_in_rsci_bdwt(ray_chan_in_rsci_bdwt),
      .ray_chan_in_rsci_bcwt(ray_chan_in_rsci_bcwt),
      .ray_chan_in_rsci_idat(ray_chan_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayOut_rsci
// ------------------------------------------------------------------


module RayCollector_run_rayOut_rsci (
  clk, arst_n, rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy, run_wen, rayOut_rsci_oswt,
      rayOut_rsci_wen_comp, rayOut_rsci_idat
);
  input clk;
  input arst_n;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;
  input run_wen;
  input rayOut_rsci_oswt;
  output rayOut_rsci_wen_comp;
  input [165:0] rayOut_rsci_idat;


  // Interconnect Declarations
  wire rayOut_rsci_irdy;
  wire rayOut_rsci_biwt;
  wire rayOut_rsci_bdwt;
  wire rayOut_rsci_bcwt;
  wire rayOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd139),
  .width(32'sd166)) rayOut_rsci (
      .irdy(rayOut_rsci_irdy),
      .ivld(rayOut_rsci_ivld_run_sct),
      .idat(rayOut_rsci_idat),
      .rdy(rayOut_rsc_rdy),
      .vld(rayOut_rsc_vld),
      .dat(rayOut_rsc_dat)
    );
  RayCollector_run_rayOut_rsci_rayOut_wait_ctrl RayCollector_run_rayOut_rsci_rayOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .rayOut_rsci_oswt(rayOut_rsci_oswt),
      .rayOut_rsci_irdy(rayOut_rsci_irdy),
      .rayOut_rsci_biwt(rayOut_rsci_biwt),
      .rayOut_rsci_bdwt(rayOut_rsci_bdwt),
      .rayOut_rsci_bcwt(rayOut_rsci_bcwt),
      .rayOut_rsci_ivld_run_sct(rayOut_rsci_ivld_run_sct)
    );
  RayCollector_run_rayOut_rsci_rayOut_wait_dp RayCollector_run_rayOut_rsci_rayOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rayOut_rsci_oswt(rayOut_rsci_oswt),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp),
      .rayOut_rsci_biwt(rayOut_rsci_biwt),
      .rayOut_rsci_bdwt(rayOut_rsci_bdwt),
      .rayOut_rsci_bcwt(rayOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsOut_rsci
// ------------------------------------------------------------------


module RayCollector_run_paramsOut_rsci (
  clk, arst_n, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy, run_wen,
      paramsOut_rsci_oswt, paramsOut_rsci_wen_comp, paramsOut_rsci_idat
);
  input clk;
  input arst_n;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  input run_wen;
  input paramsOut_rsci_oswt;
  output paramsOut_rsci_wen_comp;
  input [92:0] paramsOut_rsci_idat;


  // Interconnect Declarations
  wire paramsOut_rsci_irdy;
  wire paramsOut_rsci_biwt;
  wire paramsOut_rsci_bdwt;
  wire paramsOut_rsci_bcwt;
  wire paramsOut_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd138),
  .width(32'sd93)) paramsOut_rsci (
      .irdy(paramsOut_rsci_irdy),
      .ivld(paramsOut_rsci_ivld_run_sct),
      .idat(paramsOut_rsci_idat),
      .rdy(paramsOut_rsc_rdy),
      .vld(paramsOut_rsc_vld),
      .dat(paramsOut_rsc_dat)
    );
  RayCollector_run_paramsOut_rsci_paramsOut_wait_ctrl RayCollector_run_paramsOut_rsci_paramsOut_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_irdy(paramsOut_rsci_irdy),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt),
      .paramsOut_rsci_ivld_run_sct(paramsOut_rsci_ivld_run_sct)
    );
  RayCollector_run_paramsOut_rsci_paramsOut_wait_dp RayCollector_run_paramsOut_rsci_paramsOut_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsci_oswt(paramsOut_rsci_oswt),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_biwt(paramsOut_rsci_biwt),
      .paramsOut_rsci_bdwt(paramsOut_rsci_bdwt),
      .paramsOut_rsci_bcwt(paramsOut_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_paramsIn_rsci
// ------------------------------------------------------------------


module RayCollector_run_paramsIn_rsci (
  clk, arst_n, paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, run_wen, paramsIn_rsci_oswt,
      paramsIn_rsci_wen_comp, paramsIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [92:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  input run_wen;
  input paramsIn_rsci_oswt;
  output paramsIn_rsci_wen_comp;
  output [92:0] paramsIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire paramsIn_rsci_biwt;
  wire paramsIn_rsci_bdwt;
  wire paramsIn_rsci_bcwt;
  wire paramsIn_rsci_irdy_run_sct;
  wire paramsIn_rsci_ivld;
  wire [92:0] paramsIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd137),
  .width(32'sd93)) paramsIn_rsci (
      .rdy(paramsIn_rsc_rdy),
      .vld(paramsIn_rsc_vld),
      .dat(paramsIn_rsc_dat),
      .irdy(paramsIn_rsci_irdy_run_sct),
      .ivld(paramsIn_rsci_ivld),
      .idat(paramsIn_rsci_idat)
    );
  RayCollector_run_paramsIn_rsci_paramsIn_wait_ctrl RayCollector_run_paramsIn_rsci_paramsIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_irdy_run_sct(paramsIn_rsci_irdy_run_sct),
      .paramsIn_rsci_ivld(paramsIn_rsci_ivld)
    );
  RayCollector_run_paramsIn_rsci_paramsIn_wait_dp RayCollector_run_paramsIn_rsci_paramsIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsci_oswt(paramsIn_rsci_oswt),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt),
      .paramsIn_rsci_biwt(paramsIn_rsci_biwt),
      .paramsIn_rsci_bdwt(paramsIn_rsci_bdwt),
      .paramsIn_rsci_bcwt(paramsIn_rsci_bcwt),
      .paramsIn_rsci_idat(paramsIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run_rayIn_rsci
// ------------------------------------------------------------------


module RayCollector_run_rayIn_rsci (
  clk, arst_n, rayIn_rsc_dat, rayIn_rsc_vld, rayIn_rsc_rdy, run_wen, rayIn_rsci_oswt,
      rayIn_rsci_wen_comp, rayIn_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [165:0] rayIn_rsc_dat;
  input rayIn_rsc_vld;
  output rayIn_rsc_rdy;
  input run_wen;
  input rayIn_rsci_oswt;
  output rayIn_rsci_wen_comp;
  output [165:0] rayIn_rsci_idat_mxwt;


  // Interconnect Declarations
  wire rayIn_rsci_biwt;
  wire rayIn_rsci_bdwt;
  wire rayIn_rsci_bcwt;
  wire rayIn_rsci_irdy_run_sct;
  wire rayIn_rsci_ivld;
  wire [165:0] rayIn_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd136),
  .width(32'sd166)) rayIn_rsci (
      .rdy(rayIn_rsc_rdy),
      .vld(rayIn_rsc_vld),
      .dat(rayIn_rsc_dat),
      .irdy(rayIn_rsci_irdy_run_sct),
      .ivld(rayIn_rsci_ivld),
      .idat(rayIn_rsci_idat)
    );
  RayCollector_run_rayIn_rsci_rayIn_wait_ctrl RayCollector_run_rayIn_rsci_rayIn_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .rayIn_rsci_oswt(rayIn_rsci_oswt),
      .rayIn_rsci_biwt(rayIn_rsci_biwt),
      .rayIn_rsci_bdwt(rayIn_rsci_bdwt),
      .rayIn_rsci_bcwt(rayIn_rsci_bcwt),
      .rayIn_rsci_irdy_run_sct(rayIn_rsci_irdy_run_sct),
      .rayIn_rsci_ivld(rayIn_rsci_ivld)
    );
  RayCollector_run_rayIn_rsci_rayIn_wait_dp RayCollector_run_rayIn_rsci_rayIn_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .rayIn_rsci_oswt(rayIn_rsci_oswt),
      .rayIn_rsci_wen_comp(rayIn_rsci_wen_comp),
      .rayIn_rsci_idat_mxwt(rayIn_rsci_idat_mxwt),
      .rayIn_rsci_biwt(rayIn_rsci_biwt),
      .rayIn_rsci_bdwt(rayIn_rsci_bdwt),
      .rayIn_rsci_bcwt(rayIn_rsci_bcwt),
      .rayIn_rsci_idat(rayIn_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_output_pxl_serial_rsci
// ------------------------------------------------------------------


module PixelAccumulator_run_output_pxl_serial_rsci (
  clk, arst_n, output_pxl_serial_rsc_dat, output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy,
      run_wen, output_pxl_serial_rsci_oswt, output_pxl_serial_rsci_wen_comp, output_pxl_serial_rsci_idat
);
  input clk;
  input arst_n;
  output [23:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;
  input run_wen;
  input output_pxl_serial_rsci_oswt;
  output output_pxl_serial_rsci_wen_comp;
  input [23:0] output_pxl_serial_rsci_idat;


  // Interconnect Declarations
  wire output_pxl_serial_rsci_irdy;
  wire output_pxl_serial_rsci_biwt;
  wire output_pxl_serial_rsci_bdwt;
  wire output_pxl_serial_rsci_bcwt;
  wire output_pxl_serial_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd151),
  .width(32'sd24)) output_pxl_serial_rsci (
      .irdy(output_pxl_serial_rsci_irdy),
      .ivld(output_pxl_serial_rsci_ivld_run_sct),
      .idat(output_pxl_serial_rsci_idat),
      .rdy(output_pxl_serial_rsc_rdy),
      .vld(output_pxl_serial_rsc_vld),
      .dat(output_pxl_serial_rsc_dat)
    );
  PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .output_pxl_serial_rsci_oswt(output_pxl_serial_rsci_oswt),
      .output_pxl_serial_rsci_irdy(output_pxl_serial_rsci_irdy),
      .output_pxl_serial_rsci_biwt(output_pxl_serial_rsci_biwt),
      .output_pxl_serial_rsci_bdwt(output_pxl_serial_rsci_bdwt),
      .output_pxl_serial_rsci_bcwt(output_pxl_serial_rsci_bcwt),
      .output_pxl_serial_rsci_ivld_run_sct(output_pxl_serial_rsci_ivld_run_sct)
    );
  PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp PixelAccumulator_run_output_pxl_serial_rsci_output_pxl_serial_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_pxl_serial_rsci_oswt(output_pxl_serial_rsci_oswt),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp),
      .output_pxl_serial_rsci_biwt(output_pxl_serial_rsci_biwt),
      .output_pxl_serial_rsci_bdwt(output_pxl_serial_rsci_bdwt),
      .output_pxl_serial_rsci_bcwt(output_pxl_serial_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_pxl_sample_rsci
// ------------------------------------------------------------------


module PixelAccumulator_run_pxl_sample_rsci (
  clk, arst_n, pxl_sample_rsc_dat, pxl_sample_rsc_vld, pxl_sample_rsc_rdy, run_wen,
      pxl_sample_rsci_oswt, pxl_sample_rsci_wen_comp, pxl_sample_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [80:0] pxl_sample_rsc_dat;
  input pxl_sample_rsc_vld;
  output pxl_sample_rsc_rdy;
  input run_wen;
  input pxl_sample_rsci_oswt;
  output pxl_sample_rsci_wen_comp;
  output [80:0] pxl_sample_rsci_idat_mxwt;


  // Interconnect Declarations
  wire pxl_sample_rsci_biwt;
  wire pxl_sample_rsci_bdwt;
  wire pxl_sample_rsci_bcwt;
  wire pxl_sample_rsci_irdy_run_sct;
  wire pxl_sample_rsci_ivld;
  wire [80:0] pxl_sample_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd150),
  .width(32'sd81)) pxl_sample_rsci (
      .rdy(pxl_sample_rsc_rdy),
      .vld(pxl_sample_rsc_vld),
      .dat(pxl_sample_rsc_dat),
      .irdy(pxl_sample_rsci_irdy_run_sct),
      .ivld(pxl_sample_rsci_ivld),
      .idat(pxl_sample_rsci_idat)
    );
  PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_ctrl PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .pxl_sample_rsci_oswt(pxl_sample_rsci_oswt),
      .pxl_sample_rsci_biwt(pxl_sample_rsci_biwt),
      .pxl_sample_rsci_bdwt(pxl_sample_rsci_bdwt),
      .pxl_sample_rsci_bcwt(pxl_sample_rsci_bcwt),
      .pxl_sample_rsci_irdy_run_sct(pxl_sample_rsci_irdy_run_sct),
      .pxl_sample_rsci_ivld(pxl_sample_rsci_ivld)
    );
  PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_dp PixelAccumulator_run_pxl_sample_rsci_pxl_sample_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .pxl_sample_rsci_oswt(pxl_sample_rsci_oswt),
      .pxl_sample_rsci_wen_comp(pxl_sample_rsci_wen_comp),
      .pxl_sample_rsci_idat_mxwt(pxl_sample_rsci_idat_mxwt),
      .pxl_sample_rsci_biwt(pxl_sample_rsci_biwt),
      .pxl_sample_rsci_bdwt(pxl_sample_rsci_bdwt),
      .pxl_sample_rsci_bcwt(pxl_sample_rsci_bcwt),
      .pxl_sample_rsci_idat(pxl_sample_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run_accumulator_parms_rsci
// ------------------------------------------------------------------


module PixelAccumulator_run_accumulator_parms_rsci (
  clk, arst_n, accumulator_parms_rsc_dat, accumulator_parms_rsc_vld, accumulator_parms_rsc_rdy,
      run_wen, accumulator_parms_rsci_oswt, accumulator_parms_rsci_wen_comp, accumulator_parms_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [419:0] accumulator_parms_rsc_dat;
  input accumulator_parms_rsc_vld;
  output accumulator_parms_rsc_rdy;
  input run_wen;
  input accumulator_parms_rsci_oswt;
  output accumulator_parms_rsci_wen_comp;
  output [34:0] accumulator_parms_rsci_idat_mxwt;


  // Interconnect Declarations
  wire accumulator_parms_rsci_biwt;
  wire accumulator_parms_rsci_bdwt;
  wire accumulator_parms_rsci_bcwt;
  wire accumulator_parms_rsci_irdy_run_sct;
  wire accumulator_parms_rsci_ivld;
  wire [419:0] accumulator_parms_rsci_idat;
  wire [34:0] accumulator_parms_rsci_idat_mxwt_pconst;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd149),
  .width(32'sd420)) accumulator_parms_rsci (
      .rdy(accumulator_parms_rsc_rdy),
      .vld(accumulator_parms_rsc_vld),
      .dat(accumulator_parms_rsc_dat),
      .irdy(accumulator_parms_rsci_irdy_run_sct),
      .ivld(accumulator_parms_rsci_ivld),
      .idat(accumulator_parms_rsci_idat)
    );
  PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_ctrl PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .accumulator_parms_rsci_oswt(accumulator_parms_rsci_oswt),
      .accumulator_parms_rsci_biwt(accumulator_parms_rsci_biwt),
      .accumulator_parms_rsci_bdwt(accumulator_parms_rsci_bdwt),
      .accumulator_parms_rsci_bcwt(accumulator_parms_rsci_bcwt),
      .accumulator_parms_rsci_irdy_run_sct(accumulator_parms_rsci_irdy_run_sct),
      .accumulator_parms_rsci_ivld(accumulator_parms_rsci_ivld)
    );
  PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_dp PixelAccumulator_run_accumulator_parms_rsci_accumulator_parms_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulator_parms_rsci_oswt(accumulator_parms_rsci_oswt),
      .accumulator_parms_rsci_wen_comp(accumulator_parms_rsci_wen_comp),
      .accumulator_parms_rsci_idat_mxwt(accumulator_parms_rsci_idat_mxwt_pconst),
      .accumulator_parms_rsci_biwt(accumulator_parms_rsci_biwt),
      .accumulator_parms_rsci_bdwt(accumulator_parms_rsci_bdwt),
      .accumulator_parms_rsci_bcwt(accumulator_parms_rsci_bcwt),
      .accumulator_parms_rsci_idat(accumulator_parms_rsci_idat)
    );
  assign accumulator_parms_rsci_idat_mxwt = accumulator_parms_rsci_idat_mxwt_pconst;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer_run
// ------------------------------------------------------------------


module ParamsDeserializer_run (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      qbuffer_params_rsc_dat, qbuffer_params_rsc_vld, qbuffer_params_rsc_rdy, render_params_rsc_dat,
      render_params_rsc_vld, render_params_rsc_rdy, accum_params_rsc_dat, accum_params_rsc_vld,
      accum_params_rsc_rdy, quad_serial_out_rsc_dat, quad_serial_out_rsc_vld, quad_serial_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [11:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [56:0] qbuffer_params_rsc_dat;
  output qbuffer_params_rsc_vld;
  input qbuffer_params_rsc_rdy;
  output [419:0] render_params_rsc_dat;
  output render_params_rsc_vld;
  input render_params_rsc_rdy;
  output [419:0] accum_params_rsc_dat;
  output accum_params_rsc_vld;
  input accum_params_rsc_rdy;
  output [376:0] quad_serial_out_rsc_dat;
  output quad_serial_out_rsc_vld;
  input quad_serial_out_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire inputChannel_rsci_wen_comp;
  wire [11:0] inputChannel_rsci_idat_mxwt;
  wire qbuffer_params_rsci_wen_comp;
  wire render_params_rsci_wen_comp;
  wire accum_params_rsci_wen_comp;
  wire quad_serial_out_rsci_wen_comp;
  reg [10:0] qbuffer_params_rsci_idat_56_46;
  reg [10:0] qbuffer_params_rsci_idat_45_35;
  reg [1:0] qbuffer_params_rsci_idat_12_11;
  reg [10:0] qbuffer_params_rsci_idat_10_0;
  reg [2:0] quad_serial_out_rsci_idat_376_374;
  reg [11:0] quad_serial_out_rsci_idat_373_362;
  reg [2:0] quad_serial_out_rsci_idat_349_347;
  reg [11:0] quad_serial_out_rsci_idat_346_335;
  reg [2:0] quad_serial_out_rsci_idat_322_320;
  reg [11:0] quad_serial_out_rsci_idat_319_308;
  reg [6:0] quad_serial_out_rsci_idat_295_289;
  reg quad_serial_out_rsci_idat_264;
  reg quad_serial_out_rsci_idat_239;
  reg quad_serial_out_rsci_idat_214;
  reg [1:0] quad_serial_out_rsci_idat_189_188;
  reg [11:0] quad_serial_out_rsci_idat_175_164;
  reg [1:0] quad_serial_out_rsci_idat_163_162;
  reg [11:0] quad_serial_out_rsci_idat_149_138;
  reg [1:0] quad_serial_out_rsci_idat_137_136;
  reg [11:0] quad_serial_out_rsci_idat_123_112;
  reg quad_serial_out_rsci_idat_111;
  reg [2:0] quad_serial_out_rsci_idat_110_108;
  wire [6:0] fsm_output;
  wire or_dcpl_7;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire or_dcpl_18;
  wire mux_tmp_7;
  wire and_dcpl_26;
  wire mux_tmp_11;
  wire or_dcpl_30;
  wire or_dcpl_40;
  wire and_dcpl_61;
  wire or_dcpl_69;
  wire quad_serial_out_and_cse;
  wire accum_params_and_cse;
  wire qbuffer_params_and_cse;
  reg reg_quad_serial_out_rsci_ivld_run_psct_cse;
  reg reg_accum_params_rsci_ivld_run_psct_cse;
  reg reg_qbuffer_params_rsci_ivld_run_psct_cse;
  reg reg_inputChannel_rsci_irdy_run_psct_cse;
  reg for_slc_for_acc_6_itm;
  reg operator_33_true_operator_33_true_and_itm;
  reg [10:0] reg_accum_params_rsci_idat_10_0_cse;
  reg [1:0] reg_accum_params_rsci_idat_12_11_cse;
  reg [11:0] reg_accum_params_rsci_idat_24_13_cse;
  reg [11:0] reg_accum_params_rsci_idat_36_25_cse;
  reg [11:0] reg_accum_params_rsci_idat_51_40_cse;
  reg [11:0] reg_accum_params_rsci_idat_63_52_cse;
  reg [11:0] reg_accum_params_rsci_idat_78_67_cse;
  reg [11:0] reg_accum_params_rsci_idat_90_79_cse;
  reg [2:0] reg_accum_params_rsci_idat_93_91_cse;
  reg [10:0] reg_accum_params_rsci_idat_126_116_cse;
  reg [10:0] reg_accum_params_rsci_idat_137_127_cse;
  reg [10:0] reg_accum_params_rsci_idat_148_138_cse;
  reg [10:0] reg_accum_params_rsci_idat_159_149_cse;
  reg [10:0] reg_accum_params_rsci_idat_170_160_cse;
  reg [10:0] reg_accum_params_rsci_idat_181_171_cse;
  reg [10:0] reg_accum_params_rsci_idat_192_182_cse;
  reg [10:0] reg_accum_params_rsci_idat_203_193_cse;
  reg [10:0] reg_accum_params_rsci_idat_214_204_cse;
  reg [10:0] reg_accum_params_rsci_idat_225_215_cse;
  reg [10:0] reg_accum_params_rsci_idat_236_226_cse;
  reg [10:0] reg_accum_params_rsci_idat_247_237_cse;
  reg [10:0] reg_accum_params_rsci_idat_258_248_cse;
  reg [10:0] reg_accum_params_rsci_idat_269_259_cse;
  reg [10:0] reg_accum_params_rsci_idat_280_270_cse;
  reg [10:0] reg_accum_params_rsci_idat_291_281_cse;
  reg [2:0] reg_accum_params_rsci_idat_294_292_cse;
  reg [10:0] reg_accum_params_rsci_idat_305_295_cse;
  reg [10:0] reg_accum_params_rsci_idat_316_306_cse;
  reg [2:0] reg_accum_params_rsci_idat_319_317_cse;
  reg [10:0] reg_accum_params_rsci_idat_330_320_cse;
  reg [10:0] reg_accum_params_rsci_idat_341_331_cse;
  reg [10:0] reg_accum_params_rsci_idat_355_345_cse;
  reg [10:0] reg_accum_params_rsci_idat_366_356_cse;
  reg [10:0] reg_accum_params_rsci_idat_380_370_cse;
  reg [10:0] reg_accum_params_rsci_idat_391_381_cse;
  reg [10:0] reg_accum_params_rsci_idat_405_395_cse;
  reg [10:0] reg_accum_params_rsci_idat_416_406_cse;
  reg [2:0] reg_accum_params_rsci_idat_419_417_cse;
  reg [11:0] for_inputChannel_tmp_11_sva;
  reg [11:0] for_inputChannel_tmp_14_sva;
  reg [11:0] for_inputChannel_tmp_17_sva;
  reg [11:0] for_quad_to_sram_quad_color_r_23_12_sva;
  reg [11:0] for_quad_to_sram_quad_color_g_23_12_sva;
  reg [11:0] for_quad_to_sram_quad_color_b_23_12_sva;
  reg [2:0] for_for_slc_for_inputChannel_tmp_37_2_0_1_itm;
  reg [2:0] for_for_slc_for_inputChannel_tmp_34_2_0_1_itm;
  reg [1:0] for_for_slc_for_inputChannel_tmp_13_1_0_1_itm;
  reg for_for_slc_for_inputChannel_tmp_10_0_1_itm;
  reg [2:0] for_for_slc_for_inputChannel_tmp_9_2_0_1_itm;
  reg [10:0] inputChannel_tmp_sva_10_0;
  reg [10:0] inputChannel_tmp_40_sva_10_0;
  reg [10:0] inputChannel_tmp_42_sva_10_0;
  reg [10:0] inputChannel_tmp_43_sva_10_0;
  wire [5:0] for_i_5_0_sva_1_mx0w1;
  wire [6:0] nl_for_i_5_0_sva_1_mx0w1;
  wire [11:0] operator_11_false_acc_sdt_sva_1;
  wire [12:0] nl_operator_11_false_acc_sdt_sva_1;
  wire not_tmp_90;
  wire [10:0] mux_225_rgt;
  wire mux_tmp_160;
  reg for_quad_to_sram_corner_pt_x_sva_11;
  reg [10:0] for_quad_to_sram_corner_pt_x_sva_10_0;
  reg for_quad_to_sram_corner_pt_y_sva_11;
  reg [10:0] for_quad_to_sram_corner_pt_y_sva_10_0;
  reg for_quad_to_sram_corner_pt_z_sva_11;
  reg [10:0] for_quad_to_sram_corner_pt_z_sva_10_0;
  reg for_quad_to_sram_u_x_sva_11;
  reg [10:0] for_quad_to_sram_u_x_sva_10_0;
  reg for_quad_to_sram_u_y_sva_11;
  reg [10:0] for_quad_to_sram_u_y_sva_10_0;
  reg for_quad_to_sram_u_z_sva_11;
  reg [10:0] for_quad_to_sram_u_z_sva_10_0;
  reg for_quad_to_sram_v_x_sva_11;
  reg [10:0] for_quad_to_sram_v_x_sva_10_0;
  reg for_quad_to_sram_v_y_sva_11;
  reg [10:0] for_quad_to_sram_v_y_sva_10_0;
  reg for_quad_to_sram_v_z_sva_11;
  reg [10:0] for_quad_to_sram_v_z_sva_10_0;
  reg for_quad_to_sram_normal_x_23_12_sva_11;
  reg [10:0] for_quad_to_sram_normal_x_23_12_sva_10_0;
  reg for_quad_to_sram_normal_y_23_12_sva_11;
  reg [10:0] for_quad_to_sram_normal_y_23_12_sva_10_0;
  reg for_quad_to_sram_normal_z_23_12_sva_11;
  reg [10:0] for_quad_to_sram_normal_z_23_12_sva_10_0;
  reg for_inputChannel_tmp_20_sva_11;
  reg [10:0] for_inputChannel_tmp_20_sva_10_0;
  reg for_quad_to_sram_w_x_23_12_sva_11;
  reg [10:0] for_quad_to_sram_w_x_23_12_sva_10_0;
  reg for_inputChannel_tmp_23_sva_11;
  reg [10:0] for_inputChannel_tmp_23_sva_10_0;
  reg for_quad_to_sram_w_y_23_12_sva_11;
  reg [10:0] for_quad_to_sram_w_y_23_12_sva_10_0;
  reg for_inputChannel_tmp_26_sva_11;
  reg [10:0] for_inputChannel_tmp_26_sva_10_0;
  reg for_quad_to_sram_w_z_23_12_sva_11;
  reg [10:0] for_quad_to_sram_w_z_23_12_sva_10_0;
  reg for_inputChannel_tmp_29_sva_11;
  reg [10:0] for_inputChannel_tmp_29_sva_10_0;
  reg for_quad_to_sram_d_plane_23_12_sva_11;
  reg [10:0] for_quad_to_sram_d_plane_23_12_sva_10_0;
  reg for_inputChannel_tmp_32_sva_11;
  reg [10:0] for_inputChannel_tmp_32_sva_10_0;
  reg for_inputChannel_tmp_35_sva_11;
  reg [10:0] for_inputChannel_tmp_35_sva_10_0;
  reg for_inputChannel_tmp_38_sva_11;
  reg [10:0] for_inputChannel_tmp_38_sva_10_0;
  reg [1:0] inputChannel_tmp_4_sva_2_1;
  reg inputChannel_tmp_4_sva_0;
  reg [1:0] inputChannel_tmp_7_sva_2_1;
  reg inputChannel_tmp_7_sva_0;
  reg [3:0] inputChannel_tmp_11_sva_10_7;
  reg [6:0] inputChannel_tmp_11_sva_6_0;
  reg [4:0] inputChannel_tmp_12_sva_10_6;
  reg [5:0] inputChannel_tmp_12_sva_5_0;
  reg inputChannel_tmp_35_sva_2;
  reg [1:0] inputChannel_tmp_35_sva_1_0;
  reg inputChannel_tmp_38_sva_2;
  reg [1:0] inputChannel_tmp_38_sva_1_0;
  reg [1:0] inputChannel_tmp_41_sva_2_1;
  reg inputChannel_tmp_41_sva_0;
  reg [4:0] qbuffer_params_rsci_idat_34_30;
  reg [5:0] qbuffer_params_rsci_idat_29_24;
  reg [3:0] qbuffer_params_rsci_idat_23_20;
  reg [6:0] qbuffer_params_rsci_idat_19_13;
  reg quad_serial_out_rsci_idat_361;
  reg [10:0] quad_serial_out_rsci_idat_360_350;
  reg quad_serial_out_rsci_idat_334;
  reg [10:0] quad_serial_out_rsci_idat_333_323;
  reg quad_serial_out_rsci_idat_307;
  reg [10:0] quad_serial_out_rsci_idat_306_296;
  reg quad_serial_out_rsci_idat_288;
  reg [10:0] quad_serial_out_rsci_idat_287_277;
  reg quad_serial_out_rsci_idat_276;
  reg [10:0] quad_serial_out_rsci_idat_275_265;
  reg quad_serial_out_rsci_idat_263;
  reg [10:0] quad_serial_out_rsci_idat_262_252;
  reg quad_serial_out_rsci_idat_251;
  reg [10:0] quad_serial_out_rsci_idat_250_240;
  reg quad_serial_out_rsci_idat_238;
  reg [10:0] quad_serial_out_rsci_idat_237_227;
  reg quad_serial_out_rsci_idat_226;
  reg [10:0] quad_serial_out_rsci_idat_225_215;
  reg quad_serial_out_rsci_idat_213;
  reg [10:0] quad_serial_out_rsci_idat_212_202;
  reg quad_serial_out_rsci_idat_201;
  reg [10:0] quad_serial_out_rsci_idat_200_190;
  reg quad_serial_out_rsci_idat_187;
  reg [10:0] quad_serial_out_rsci_idat_186_176;
  reg quad_serial_out_rsci_idat_161;
  reg [10:0] quad_serial_out_rsci_idat_160_150;
  reg quad_serial_out_rsci_idat_135;
  reg [10:0] quad_serial_out_rsci_idat_134_124;
  reg quad_serial_out_rsci_idat_107;
  reg [10:0] quad_serial_out_rsci_idat_106_96;
  reg quad_serial_out_rsci_idat_95;
  reg [10:0] quad_serial_out_rsci_idat_94_84;
  reg quad_serial_out_rsci_idat_83;
  reg [10:0] quad_serial_out_rsci_idat_82_72;
  reg quad_serial_out_rsci_idat_71;
  reg [10:0] quad_serial_out_rsci_idat_70_60;
  reg quad_serial_out_rsci_idat_59;
  reg [10:0] quad_serial_out_rsci_idat_58_48;
  reg quad_serial_out_rsci_idat_47;
  reg [10:0] quad_serial_out_rsci_idat_46_36;
  reg quad_serial_out_rsci_idat_35;
  reg [10:0] quad_serial_out_rsci_idat_34_24;
  reg quad_serial_out_rsci_idat_23;
  reg [10:0] quad_serial_out_rsci_idat_22_12;
  reg quad_serial_out_rsci_idat_11;
  reg [10:0] quad_serial_out_rsci_idat_10_0;
  reg [1:0] reg_accum_params_rsci_idat_39_37_cse_2_1;
  reg reg_accum_params_rsci_idat_39_37_cse_0;
  reg [1:0] reg_accum_params_rsci_idat_66_64_cse_2_1;
  reg reg_accum_params_rsci_idat_66_64_cse_0;
  reg [3:0] reg_accum_params_rsci_idat_104_94_cse_10_7;
  reg [6:0] reg_accum_params_rsci_idat_104_94_cse_6_0;
  reg [4:0] reg_accum_params_rsci_idat_115_105_cse_10_6;
  reg [5:0] reg_accum_params_rsci_idat_115_105_cse_5_0;
  reg reg_accum_params_rsci_idat_344_342_cse_2;
  reg [1:0] reg_accum_params_rsci_idat_344_342_cse_1_0;
  reg reg_accum_params_rsci_idat_369_367_cse_2;
  reg [1:0] reg_accum_params_rsci_idat_369_367_cse_1_0;
  reg [1:0] reg_accum_params_rsci_idat_394_392_cse_2_1;
  reg reg_accum_params_rsci_idat_394_392_cse_0;
  wire nor_168_cse;
  wire nand_52_cse;
  wire and_383_cse;
  wire or_338_cse;
  wire or_216_cse;
  wire or_214_cse;
  wire nor_177_cse;
  wire and_369_cse;
  wire or_42_cse;
  wire nor_164_cse;
  wire nor_148_cse;
  wire or_178_cse;
  wire and_377_cse;
  wire and_380_cse;
  wire xnor_2_cse;
  wire or_326_cse;
  wire nor_138_cse;
  wire and_354_cse;
  wire or_285_cse;
  wire nand_53_cse;
  wire nor_125_cse;
  wire nand_44_cse;
  wire nand_33_cse;
  wire nor_173_cse;
  wire and_356_cse;
  wire or_314_cse;
  wire and_348_cse;
  wire and_131_cse;
  wire mux_248_cse;
  wire or_311_cse;
  wire mux_272_cse;
  wire and_372_cse;
  wire mux_290_cse;
  wire nand_38_cse;
  wire nor_149_cse;

  wire[0:0] mux_117_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] or_23_nl;
  wire[0:0] mux_115_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] or_31_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] or_36_nl;
  wire[0:0] or_35_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] or_169_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_27_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] or_48_nl;
  wire[0:0] or_47_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] or_51_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] or_173_nl;
  wire[0:0] or_172_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] or_171_nl;
  wire[0:0] or_170_nl;
  wire[0:0] and_31_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] or_339_nl;
  wire[0:0] nand_54_nl;
  wire[0:0] mux_132_nl;
  wire[0:0] or_57_nl;
  wire[0:0] or_56_nl;
  wire[0:0] mux_133_nl;
  wire[0:0] or_66_nl;
  wire[0:0] or_65_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] nor_174_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] and_382_nl;
  wire[0:0] nor_175_nl;
  wire[5:0] for_i_for_i_and_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] and_135_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] and_132_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] or_179_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] nor_172_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] and_378_nl;
  wire[0:0] or_182_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] nor_170_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] or_337_nl;
  wire[0:0] nor_169_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] and_376_nl;
  wire[0:0] nor_167_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] nor_166_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] nor_162_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] and_374_nl;
  wire[0:0] nor_161_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] nor_157_nl;
  wire[0:0] nor_158_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] and_373_nl;
  wire[0:0] nor_156_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] nor_153_nl;
  wire[0:0] nor_154_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] or_215_nl;
  wire[0:0] or_212_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] or_218_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] and_368_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_62_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_150_nl;
  wire[0:0] nor_151_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] and_365_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] nand_46_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] and_361_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] and_359_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] nor_140_nl;
  wire[0:0] nor_141_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] and_357_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] nand_42_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] or_248_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] nand_40_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_252_nl;
  wire[0:0] or_250_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] and_353_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] nor_137_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] nor_135_nl;
  wire[0:0] nor_136_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] and_385_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] nor_133_nl;
  wire[0:0] nor_134_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] nor_130_nl;
  wire[0:0] nor_131_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] and_349_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] nor_129_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] nor_128_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] nor_127_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] or_127_nl;
  wire[0:0] or_126_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] nand_34_nl;
  wire[0:0] nor_124_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] and_346_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] and_344_nl;
  wire[0:0] nor_122_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] or_313_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] or_282_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] and_342_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_119_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] or_308_nl;
  wire[0:0] or_309_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] nor_115_nl;
  wire[0:0] nor_116_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] nor_117_nl;
  wire[0:0] and_341_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] and_340_nl;
  wire[0:0] nor_114_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] and_339_nl;
  wire[0:0] nor_113_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] or_305_nl;
  wire[0:0] or_306_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_110_nl;
  wire[0:0] nor_111_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] nand_28_nl;
  wire[0:0] and_111_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] or_304_nl;
  wire[6:0] for_acc_nl;
  wire[7:0] nl_for_acc_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] or_155_nl;
  wire[0:0] or_26_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] or_25_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [56:0] nl_ParamsDeserializer_run_qbuffer_params_rsci_inst_qbuffer_params_rsci_idat;
  assign nl_ParamsDeserializer_run_qbuffer_params_rsci_inst_qbuffer_params_rsci_idat
      = {qbuffer_params_rsci_idat_56_46 , qbuffer_params_rsci_idat_45_35 , qbuffer_params_rsci_idat_34_30
      , qbuffer_params_rsci_idat_29_24 , qbuffer_params_rsci_idat_23_20 , qbuffer_params_rsci_idat_19_13
      , qbuffer_params_rsci_idat_12_11 , qbuffer_params_rsci_idat_10_0};
  wire [419:0] nl_ParamsDeserializer_run_render_params_rsci_inst_render_params_rsci_idat;
  assign nl_ParamsDeserializer_run_render_params_rsci_inst_render_params_rsci_idat
      = {reg_accum_params_rsci_idat_419_417_cse , reg_accum_params_rsci_idat_416_406_cse
      , reg_accum_params_rsci_idat_405_395_cse , reg_accum_params_rsci_idat_394_392_cse_2_1
      , reg_accum_params_rsci_idat_394_392_cse_0 , reg_accum_params_rsci_idat_391_381_cse
      , reg_accum_params_rsci_idat_380_370_cse , reg_accum_params_rsci_idat_369_367_cse_2
      , reg_accum_params_rsci_idat_369_367_cse_1_0 , reg_accum_params_rsci_idat_366_356_cse
      , reg_accum_params_rsci_idat_355_345_cse , reg_accum_params_rsci_idat_344_342_cse_2
      , reg_accum_params_rsci_idat_344_342_cse_1_0 , reg_accum_params_rsci_idat_341_331_cse
      , reg_accum_params_rsci_idat_330_320_cse , reg_accum_params_rsci_idat_319_317_cse
      , reg_accum_params_rsci_idat_316_306_cse , reg_accum_params_rsci_idat_305_295_cse
      , reg_accum_params_rsci_idat_294_292_cse , reg_accum_params_rsci_idat_291_281_cse
      , reg_accum_params_rsci_idat_280_270_cse , reg_accum_params_rsci_idat_269_259_cse
      , reg_accum_params_rsci_idat_258_248_cse , reg_accum_params_rsci_idat_247_237_cse
      , reg_accum_params_rsci_idat_236_226_cse , reg_accum_params_rsci_idat_225_215_cse
      , reg_accum_params_rsci_idat_214_204_cse , reg_accum_params_rsci_idat_203_193_cse
      , reg_accum_params_rsci_idat_192_182_cse , reg_accum_params_rsci_idat_181_171_cse
      , reg_accum_params_rsci_idat_170_160_cse , reg_accum_params_rsci_idat_159_149_cse
      , reg_accum_params_rsci_idat_148_138_cse , reg_accum_params_rsci_idat_137_127_cse
      , reg_accum_params_rsci_idat_126_116_cse , reg_accum_params_rsci_idat_115_105_cse_10_6
      , reg_accum_params_rsci_idat_115_105_cse_5_0 , reg_accum_params_rsci_idat_104_94_cse_10_7
      , reg_accum_params_rsci_idat_104_94_cse_6_0 , reg_accum_params_rsci_idat_93_91_cse
      , reg_accum_params_rsci_idat_90_79_cse , reg_accum_params_rsci_idat_78_67_cse
      , reg_accum_params_rsci_idat_66_64_cse_2_1 , reg_accum_params_rsci_idat_66_64_cse_0
      , reg_accum_params_rsci_idat_63_52_cse , reg_accum_params_rsci_idat_51_40_cse
      , reg_accum_params_rsci_idat_39_37_cse_2_1 , reg_accum_params_rsci_idat_39_37_cse_0
      , reg_accum_params_rsci_idat_36_25_cse , reg_accum_params_rsci_idat_24_13_cse
      , reg_accum_params_rsci_idat_12_11_cse , reg_accum_params_rsci_idat_10_0_cse};
  wire [419:0] nl_ParamsDeserializer_run_accum_params_rsci_inst_accum_params_rsci_idat;
  assign nl_ParamsDeserializer_run_accum_params_rsci_inst_accum_params_rsci_idat
      = {reg_accum_params_rsci_idat_419_417_cse , reg_accum_params_rsci_idat_416_406_cse
      , reg_accum_params_rsci_idat_405_395_cse , reg_accum_params_rsci_idat_394_392_cse_2_1
      , reg_accum_params_rsci_idat_394_392_cse_0 , reg_accum_params_rsci_idat_391_381_cse
      , reg_accum_params_rsci_idat_380_370_cse , reg_accum_params_rsci_idat_369_367_cse_2
      , reg_accum_params_rsci_idat_369_367_cse_1_0 , reg_accum_params_rsci_idat_366_356_cse
      , reg_accum_params_rsci_idat_355_345_cse , reg_accum_params_rsci_idat_344_342_cse_2
      , reg_accum_params_rsci_idat_344_342_cse_1_0 , reg_accum_params_rsci_idat_341_331_cse
      , reg_accum_params_rsci_idat_330_320_cse , reg_accum_params_rsci_idat_319_317_cse
      , reg_accum_params_rsci_idat_316_306_cse , reg_accum_params_rsci_idat_305_295_cse
      , reg_accum_params_rsci_idat_294_292_cse , reg_accum_params_rsci_idat_291_281_cse
      , reg_accum_params_rsci_idat_280_270_cse , reg_accum_params_rsci_idat_269_259_cse
      , reg_accum_params_rsci_idat_258_248_cse , reg_accum_params_rsci_idat_247_237_cse
      , reg_accum_params_rsci_idat_236_226_cse , reg_accum_params_rsci_idat_225_215_cse
      , reg_accum_params_rsci_idat_214_204_cse , reg_accum_params_rsci_idat_203_193_cse
      , reg_accum_params_rsci_idat_192_182_cse , reg_accum_params_rsci_idat_181_171_cse
      , reg_accum_params_rsci_idat_170_160_cse , reg_accum_params_rsci_idat_159_149_cse
      , reg_accum_params_rsci_idat_148_138_cse , reg_accum_params_rsci_idat_137_127_cse
      , reg_accum_params_rsci_idat_126_116_cse , reg_accum_params_rsci_idat_115_105_cse_10_6
      , reg_accum_params_rsci_idat_115_105_cse_5_0 , reg_accum_params_rsci_idat_104_94_cse_10_7
      , reg_accum_params_rsci_idat_104_94_cse_6_0 , reg_accum_params_rsci_idat_93_91_cse
      , reg_accum_params_rsci_idat_90_79_cse , reg_accum_params_rsci_idat_78_67_cse
      , reg_accum_params_rsci_idat_66_64_cse_2_1 , reg_accum_params_rsci_idat_66_64_cse_0
      , reg_accum_params_rsci_idat_63_52_cse , reg_accum_params_rsci_idat_51_40_cse
      , reg_accum_params_rsci_idat_39_37_cse_2_1 , reg_accum_params_rsci_idat_39_37_cse_0
      , reg_accum_params_rsci_idat_36_25_cse , reg_accum_params_rsci_idat_24_13_cse
      , reg_accum_params_rsci_idat_12_11_cse , reg_accum_params_rsci_idat_10_0_cse};
  wire [376:0] nl_ParamsDeserializer_run_quad_serial_out_rsci_inst_quad_serial_out_rsci_idat;
  assign nl_ParamsDeserializer_run_quad_serial_out_rsci_inst_quad_serial_out_rsci_idat
      = {quad_serial_out_rsci_idat_376_374 , quad_serial_out_rsci_idat_373_362 ,
      quad_serial_out_rsci_idat_361 , quad_serial_out_rsci_idat_360_350 , quad_serial_out_rsci_idat_349_347
      , quad_serial_out_rsci_idat_346_335 , quad_serial_out_rsci_idat_334 , quad_serial_out_rsci_idat_333_323
      , quad_serial_out_rsci_idat_322_320 , quad_serial_out_rsci_idat_319_308 , quad_serial_out_rsci_idat_307
      , quad_serial_out_rsci_idat_306_296 , quad_serial_out_rsci_idat_295_289 , quad_serial_out_rsci_idat_288
      , quad_serial_out_rsci_idat_287_277 , quad_serial_out_rsci_idat_276 , quad_serial_out_rsci_idat_275_265
      , quad_serial_out_rsci_idat_264 , quad_serial_out_rsci_idat_263 , quad_serial_out_rsci_idat_262_252
      , quad_serial_out_rsci_idat_251 , quad_serial_out_rsci_idat_250_240 , quad_serial_out_rsci_idat_239
      , quad_serial_out_rsci_idat_238 , quad_serial_out_rsci_idat_237_227 , quad_serial_out_rsci_idat_226
      , quad_serial_out_rsci_idat_225_215 , quad_serial_out_rsci_idat_214 , quad_serial_out_rsci_idat_213
      , quad_serial_out_rsci_idat_212_202 , quad_serial_out_rsci_idat_201 , quad_serial_out_rsci_idat_200_190
      , quad_serial_out_rsci_idat_189_188 , quad_serial_out_rsci_idat_187 , quad_serial_out_rsci_idat_186_176
      , quad_serial_out_rsci_idat_175_164 , quad_serial_out_rsci_idat_163_162 , quad_serial_out_rsci_idat_161
      , quad_serial_out_rsci_idat_160_150 , quad_serial_out_rsci_idat_149_138 , quad_serial_out_rsci_idat_137_136
      , quad_serial_out_rsci_idat_135 , quad_serial_out_rsci_idat_134_124 , quad_serial_out_rsci_idat_123_112
      , quad_serial_out_rsci_idat_111 , quad_serial_out_rsci_idat_110_108 , quad_serial_out_rsci_idat_107
      , quad_serial_out_rsci_idat_106_96 , quad_serial_out_rsci_idat_95 , quad_serial_out_rsci_idat_94_84
      , quad_serial_out_rsci_idat_83 , quad_serial_out_rsci_idat_82_72 , quad_serial_out_rsci_idat_71
      , quad_serial_out_rsci_idat_70_60 , quad_serial_out_rsci_idat_59 , quad_serial_out_rsci_idat_58_48
      , quad_serial_out_rsci_idat_47 , quad_serial_out_rsci_idat_46_36 , quad_serial_out_rsci_idat_35
      , quad_serial_out_rsci_idat_34_24 , quad_serial_out_rsci_idat_23 , quad_serial_out_rsci_idat_22_12
      , quad_serial_out_rsci_idat_11 , quad_serial_out_rsci_idat_10_0};
  wire [0:0] nl_ParamsDeserializer_run_run_fsm_inst_for_C_41_tr0;
  assign nl_ParamsDeserializer_run_run_fsm_inst_for_C_41_tr0 = operator_33_true_operator_33_true_and_itm
      | (~ for_slc_for_acc_6_itm);
  ParamsDeserializer_run_inputChannel_rsci ParamsDeserializer_run_inputChannel_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .run_wen(run_wen),
      .inputChannel_rsci_oswt(reg_inputChannel_rsci_irdy_run_psct_cse),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .inputChannel_rsci_idat_mxwt(inputChannel_rsci_idat_mxwt)
    );
  ParamsDeserializer_run_qbuffer_params_rsci ParamsDeserializer_run_qbuffer_params_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .qbuffer_params_rsc_dat(qbuffer_params_rsc_dat),
      .qbuffer_params_rsc_vld(qbuffer_params_rsc_vld),
      .qbuffer_params_rsc_rdy(qbuffer_params_rsc_rdy),
      .run_wen(run_wen),
      .qbuffer_params_rsci_oswt(reg_qbuffer_params_rsci_ivld_run_psct_cse),
      .qbuffer_params_rsci_wen_comp(qbuffer_params_rsci_wen_comp),
      .qbuffer_params_rsci_idat(nl_ParamsDeserializer_run_qbuffer_params_rsci_inst_qbuffer_params_rsci_idat[56:0])
    );
  ParamsDeserializer_run_render_params_rsci ParamsDeserializer_run_render_params_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsc_dat(render_params_rsc_dat),
      .render_params_rsc_vld(render_params_rsc_vld),
      .render_params_rsc_rdy(render_params_rsc_rdy),
      .run_wen(run_wen),
      .render_params_rsci_oswt(reg_accum_params_rsci_ivld_run_psct_cse),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .render_params_rsci_idat(nl_ParamsDeserializer_run_render_params_rsci_inst_render_params_rsci_idat[419:0])
    );
  ParamsDeserializer_run_accum_params_rsci ParamsDeserializer_run_accum_params_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accum_params_rsc_dat(accum_params_rsc_dat),
      .accum_params_rsc_vld(accum_params_rsc_vld),
      .accum_params_rsc_rdy(accum_params_rsc_rdy),
      .run_wen(run_wen),
      .accum_params_rsci_oswt(reg_accum_params_rsci_ivld_run_psct_cse),
      .accum_params_rsci_wen_comp(accum_params_rsci_wen_comp),
      .accum_params_rsci_idat(nl_ParamsDeserializer_run_accum_params_rsci_inst_accum_params_rsci_idat[419:0])
    );
  ParamsDeserializer_run_quad_serial_out_rsci ParamsDeserializer_run_quad_serial_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_serial_out_rsc_dat(quad_serial_out_rsc_dat),
      .quad_serial_out_rsc_vld(quad_serial_out_rsc_vld),
      .quad_serial_out_rsc_rdy(quad_serial_out_rsc_rdy),
      .run_wen(run_wen),
      .quad_serial_out_rsci_oswt(reg_quad_serial_out_rsci_ivld_run_psct_cse),
      .quad_serial_out_rsci_wen_comp(quad_serial_out_rsci_wen_comp),
      .quad_serial_out_rsci_idat(nl_ParamsDeserializer_run_quad_serial_out_rsci_inst_quad_serial_out_rsci_idat[376:0])
    );
  ParamsDeserializer_run_staller ParamsDeserializer_run_staller_inst (
      .run_wen(run_wen),
      .inputChannel_rsci_wen_comp(inputChannel_rsci_wen_comp),
      .qbuffer_params_rsci_wen_comp(qbuffer_params_rsci_wen_comp),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .accum_params_rsci_wen_comp(accum_params_rsci_wen_comp),
      .quad_serial_out_rsci_wen_comp(quad_serial_out_rsci_wen_comp)
    );
  ParamsDeserializer_run_run_fsm ParamsDeserializer_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_41_tr0(nl_ParamsDeserializer_run_run_fsm_inst_for_C_41_tr0[0:0])
    );
  assign quad_serial_out_and_cse = run_wen & (~(or_dcpl_7 | nand_44_cse | or_214_cse
      | (~ (fsm_output[6]))));
  assign accum_params_and_cse = run_wen & (~(or_dcpl_12 | nand_44_cse | or_dcpl_11));
  assign qbuffer_params_and_cse = run_wen & (~(or_dcpl_18 | (fsm_output[6:4]!=3'b000)));
  assign or_42_cse = (fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]);
  assign nor_177_cse = ~((fsm_output[3]) | (fsm_output[1]));
  assign and_383_cse = (fsm_output[1:0]==2'b11);
  assign and_131_cse = (fsm_output[3:1]==3'b111);
  assign nand_53_cse = ~((fsm_output[2:0]==3'b111));
  assign nor_173_cse = ~((fsm_output[5:4]!=2'b00));
  assign and_135_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[0]) & (fsm_output[3])
      & (fsm_output[1]);
  assign mux_215_nl = MUX_s_1_2_2((and_135_nl), (fsm_output[5]), fsm_output[4]);
  assign mux_216_nl = MUX_s_1_2_2((mux_215_nl), (~ mux_tmp_7), fsm_output[6]);
  assign for_i_for_i_and_nl = MUX_v_6_2_2(6'b000000, for_i_5_0_sva_1_mx0w1, (mux_216_nl));
  assign and_132_nl = (fsm_output[5]) & (fsm_output[2]) & (fsm_output[3]) & (fsm_output[1]);
  assign mux_136_nl = MUX_s_1_2_2((and_132_nl), (fsm_output[5]), fsm_output[4]);
  assign mux_137_nl = MUX_s_1_2_2((mux_136_nl), (~ mux_tmp_7), fsm_output[6]);
  assign mux_225_rgt = MUX_v_11_2_2((inputChannel_rsci_idat_mxwt[10:0]), ({5'b00000
      , (for_i_for_i_and_nl)}), mux_137_nl);
  assign or_178_cse = (fsm_output[2:0]!=3'b000);
  assign and_380_cse = (fsm_output[0]) & (fsm_output[2]);
  assign mux_248_cse = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[5]);
  assign nand_52_cse = ~((fsm_output[3:2]==2'b11));
  assign or_338_cse = (fsm_output[1:0]!=2'b00);
  assign nor_168_cse = ~((fsm_output[4]) | ((fsm_output[3]) & or_338_cse & (fsm_output[2])));
  assign and_377_cse = (fsm_output[3:0]==4'b1111);
  assign nor_164_cse = ~((fsm_output[2:1]!=2'b00));
  assign or_216_cse = (fsm_output[5:4]!=2'b10);
  assign or_214_cse = (fsm_output[5:4]!=2'b01);
  assign and_372_cse = or_338_cse & (fsm_output[3]);
  assign mux_272_cse = MUX_s_1_2_2(mux_248_cse, or_214_cse, and_372_cse);
  assign and_369_cse = (fsm_output[2:1]==2'b11);
  assign nor_149_cse = ~(and_372_cse | (fsm_output[4]));
  assign nor_148_cse = ~((fsm_output[6]) | (fsm_output[3]));
  assign mux_290_cse = MUX_s_1_2_2(and_369_cse, nor_164_cse, fsm_output[5]);
  assign or_326_cse = ((fsm_output[2:0]==3'b111)) | (fsm_output[3]);
  assign nand_44_cse = ~((fsm_output[2]) & (fsm_output[0]));
  assign and_356_cse = (fsm_output[1]) & (fsm_output[3]);
  assign nor_138_cse = ~((fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]));
  assign and_354_cse = (fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]);
  assign nand_38_cse = ~(or_338_cse & (fsm_output[3:2]==2'b11));
  assign and_348_cse = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]);
  assign nor_125_cse = ~((fsm_output[2]) | (fsm_output[0]));
  assign or_314_cse = (fsm_output[1]) | (fsm_output[3]);
  assign xnor_2_cse = ~((fsm_output[2]) ^ (fsm_output[4]));
  assign nand_33_cse = ~((fsm_output[1]) & (fsm_output[3]));
  assign or_285_cse = (fsm_output[6:5]!=2'b10);
  assign or_311_cse = (fsm_output[6:5]!=2'b01);
  assign nl_for_i_5_0_sva_1_mx0w1 = inputChannel_tmp_12_sva_5_0 + 6'b000001;
  assign for_i_5_0_sva_1_mx0w1 = nl_for_i_5_0_sva_1_mx0w1[5:0];
  assign nl_operator_11_false_acc_sdt_sva_1 = conv_u2s_11_12(inputChannel_tmp_sva_10_0)
      + 12'b111111111111;
  assign operator_11_false_acc_sdt_sva_1 = nl_operator_11_false_acc_sdt_sva_1[11:0];
  assign or_dcpl_7 = (~ (fsm_output[1])) | (fsm_output[3]);
  assign or_dcpl_11 = (fsm_output[6:4]!=3'b010);
  assign or_dcpl_12 = (fsm_output[1]) | (~ (fsm_output[3]));
  assign or_dcpl_18 = nand_33_cse | nand_44_cse;
  assign or_25_nl = (fsm_output[2]) | (fsm_output[0]);
  assign mux_118_nl = MUX_s_1_2_2(and_356_cse, (fsm_output[3]), or_25_nl);
  assign or_26_nl = (fsm_output[5]) | (mux_118_nl);
  assign mux_tmp_7 = MUX_s_1_2_2((fsm_output[5]), (or_26_nl), fsm_output[4]);
  assign and_dcpl_26 = (fsm_output[6:5]==2'b10);
  assign mux_tmp_11 = MUX_s_1_2_2((fsm_output[3]), or_314_cse, and_380_cse);
  assign or_dcpl_30 = or_dcpl_7 | (fsm_output[5]);
  assign or_dcpl_40 = (~ (fsm_output[0])) | (fsm_output[2]);
  assign and_dcpl_61 = (fsm_output[5:4]==2'b11);
  assign or_dcpl_69 = or_dcpl_12 | or_dcpl_40;
  assign not_tmp_90 = ~((fsm_output[6]) & (fsm_output[4]));
  assign mux_tmp_160 = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[4]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_serial_out_rsci_idat_11 <= 1'b0;
      quad_serial_out_rsci_idat_10_0 <= 11'b00000000000;
      quad_serial_out_rsci_idat_23 <= 1'b0;
      quad_serial_out_rsci_idat_22_12 <= 11'b00000000000;
      quad_serial_out_rsci_idat_35 <= 1'b0;
      quad_serial_out_rsci_idat_34_24 <= 11'b00000000000;
      quad_serial_out_rsci_idat_47 <= 1'b0;
      quad_serial_out_rsci_idat_46_36 <= 11'b00000000000;
      quad_serial_out_rsci_idat_59 <= 1'b0;
      quad_serial_out_rsci_idat_58_48 <= 11'b00000000000;
      quad_serial_out_rsci_idat_71 <= 1'b0;
      quad_serial_out_rsci_idat_70_60 <= 11'b00000000000;
      quad_serial_out_rsci_idat_83 <= 1'b0;
      quad_serial_out_rsci_idat_82_72 <= 11'b00000000000;
      quad_serial_out_rsci_idat_95 <= 1'b0;
      quad_serial_out_rsci_idat_94_84 <= 11'b00000000000;
      quad_serial_out_rsci_idat_107 <= 1'b0;
      quad_serial_out_rsci_idat_106_96 <= 11'b00000000000;
      quad_serial_out_rsci_idat_110_108 <= 3'b000;
      quad_serial_out_rsci_idat_111 <= 1'b0;
      quad_serial_out_rsci_idat_123_112 <= 12'b000000000000;
      quad_serial_out_rsci_idat_135 <= 1'b0;
      quad_serial_out_rsci_idat_134_124 <= 11'b00000000000;
      quad_serial_out_rsci_idat_137_136 <= 2'b00;
      quad_serial_out_rsci_idat_149_138 <= 12'b000000000000;
      quad_serial_out_rsci_idat_161 <= 1'b0;
      quad_serial_out_rsci_idat_160_150 <= 11'b00000000000;
      quad_serial_out_rsci_idat_163_162 <= 2'b00;
      quad_serial_out_rsci_idat_175_164 <= 12'b000000000000;
      quad_serial_out_rsci_idat_187 <= 1'b0;
      quad_serial_out_rsci_idat_186_176 <= 11'b00000000000;
      quad_serial_out_rsci_idat_189_188 <= 2'b00;
      quad_serial_out_rsci_idat_201 <= 1'b0;
      quad_serial_out_rsci_idat_200_190 <= 11'b00000000000;
      quad_serial_out_rsci_idat_213 <= 1'b0;
      quad_serial_out_rsci_idat_212_202 <= 11'b00000000000;
      quad_serial_out_rsci_idat_214 <= 1'b0;
      quad_serial_out_rsci_idat_226 <= 1'b0;
      quad_serial_out_rsci_idat_225_215 <= 11'b00000000000;
      quad_serial_out_rsci_idat_238 <= 1'b0;
      quad_serial_out_rsci_idat_237_227 <= 11'b00000000000;
      quad_serial_out_rsci_idat_239 <= 1'b0;
      quad_serial_out_rsci_idat_251 <= 1'b0;
      quad_serial_out_rsci_idat_250_240 <= 11'b00000000000;
      quad_serial_out_rsci_idat_263 <= 1'b0;
      quad_serial_out_rsci_idat_262_252 <= 11'b00000000000;
      quad_serial_out_rsci_idat_264 <= 1'b0;
      quad_serial_out_rsci_idat_276 <= 1'b0;
      quad_serial_out_rsci_idat_275_265 <= 11'b00000000000;
      quad_serial_out_rsci_idat_288 <= 1'b0;
      quad_serial_out_rsci_idat_287_277 <= 11'b00000000000;
      quad_serial_out_rsci_idat_295_289 <= 7'b0000000;
      quad_serial_out_rsci_idat_307 <= 1'b0;
      quad_serial_out_rsci_idat_306_296 <= 11'b00000000000;
      quad_serial_out_rsci_idat_319_308 <= 12'b000000000000;
      quad_serial_out_rsci_idat_322_320 <= 3'b000;
      quad_serial_out_rsci_idat_334 <= 1'b0;
      quad_serial_out_rsci_idat_333_323 <= 11'b00000000000;
      quad_serial_out_rsci_idat_346_335 <= 12'b000000000000;
      quad_serial_out_rsci_idat_349_347 <= 3'b000;
      quad_serial_out_rsci_idat_361 <= 1'b0;
      quad_serial_out_rsci_idat_360_350 <= 11'b00000000000;
      quad_serial_out_rsci_idat_373_362 <= 12'b000000000000;
      quad_serial_out_rsci_idat_376_374 <= 3'b000;
    end
    else if ( quad_serial_out_and_cse ) begin
      quad_serial_out_rsci_idat_11 <= for_quad_to_sram_corner_pt_x_sva_11;
      quad_serial_out_rsci_idat_10_0 <= for_quad_to_sram_corner_pt_x_sva_10_0;
      quad_serial_out_rsci_idat_23 <= for_quad_to_sram_corner_pt_y_sva_11;
      quad_serial_out_rsci_idat_22_12 <= for_quad_to_sram_corner_pt_y_sva_10_0;
      quad_serial_out_rsci_idat_35 <= for_quad_to_sram_corner_pt_z_sva_11;
      quad_serial_out_rsci_idat_34_24 <= for_quad_to_sram_corner_pt_z_sva_10_0;
      quad_serial_out_rsci_idat_47 <= for_quad_to_sram_u_x_sva_11;
      quad_serial_out_rsci_idat_46_36 <= for_quad_to_sram_u_x_sva_10_0;
      quad_serial_out_rsci_idat_59 <= for_quad_to_sram_u_y_sva_11;
      quad_serial_out_rsci_idat_58_48 <= for_quad_to_sram_u_y_sva_10_0;
      quad_serial_out_rsci_idat_71 <= for_quad_to_sram_u_z_sva_11;
      quad_serial_out_rsci_idat_70_60 <= for_quad_to_sram_u_z_sva_10_0;
      quad_serial_out_rsci_idat_83 <= for_quad_to_sram_v_x_sva_11;
      quad_serial_out_rsci_idat_82_72 <= for_quad_to_sram_v_x_sva_10_0;
      quad_serial_out_rsci_idat_95 <= for_quad_to_sram_v_y_sva_11;
      quad_serial_out_rsci_idat_94_84 <= for_quad_to_sram_v_y_sva_10_0;
      quad_serial_out_rsci_idat_107 <= for_quad_to_sram_v_z_sva_11;
      quad_serial_out_rsci_idat_106_96 <= for_quad_to_sram_v_z_sva_10_0;
      quad_serial_out_rsci_idat_110_108 <= for_for_slc_for_inputChannel_tmp_9_2_0_1_itm;
      quad_serial_out_rsci_idat_111 <= for_for_slc_for_inputChannel_tmp_10_0_1_itm;
      quad_serial_out_rsci_idat_123_112 <= for_inputChannel_tmp_11_sva;
      quad_serial_out_rsci_idat_135 <= for_quad_to_sram_normal_x_23_12_sva_11;
      quad_serial_out_rsci_idat_134_124 <= for_quad_to_sram_normal_x_23_12_sva_10_0;
      quad_serial_out_rsci_idat_137_136 <= for_for_slc_for_inputChannel_tmp_13_1_0_1_itm;
      quad_serial_out_rsci_idat_149_138 <= for_inputChannel_tmp_14_sva;
      quad_serial_out_rsci_idat_161 <= for_quad_to_sram_normal_y_23_12_sva_11;
      quad_serial_out_rsci_idat_160_150 <= for_quad_to_sram_normal_y_23_12_sva_10_0;
      quad_serial_out_rsci_idat_163_162 <= inputChannel_tmp_35_sva_1_0;
      quad_serial_out_rsci_idat_175_164 <= for_inputChannel_tmp_17_sva;
      quad_serial_out_rsci_idat_187 <= for_quad_to_sram_normal_z_23_12_sva_11;
      quad_serial_out_rsci_idat_186_176 <= for_quad_to_sram_normal_z_23_12_sva_10_0;
      quad_serial_out_rsci_idat_189_188 <= inputChannel_tmp_38_sva_1_0;
      quad_serial_out_rsci_idat_201 <= for_inputChannel_tmp_20_sva_11;
      quad_serial_out_rsci_idat_200_190 <= for_inputChannel_tmp_20_sva_10_0;
      quad_serial_out_rsci_idat_213 <= for_quad_to_sram_w_x_23_12_sva_11;
      quad_serial_out_rsci_idat_212_202 <= for_quad_to_sram_w_x_23_12_sva_10_0;
      quad_serial_out_rsci_idat_214 <= inputChannel_tmp_4_sva_0;
      quad_serial_out_rsci_idat_226 <= for_inputChannel_tmp_23_sva_11;
      quad_serial_out_rsci_idat_225_215 <= for_inputChannel_tmp_23_sva_10_0;
      quad_serial_out_rsci_idat_238 <= for_quad_to_sram_w_y_23_12_sva_11;
      quad_serial_out_rsci_idat_237_227 <= for_quad_to_sram_w_y_23_12_sva_10_0;
      quad_serial_out_rsci_idat_239 <= inputChannel_tmp_41_sva_0;
      quad_serial_out_rsci_idat_251 <= for_inputChannel_tmp_26_sva_11;
      quad_serial_out_rsci_idat_250_240 <= for_inputChannel_tmp_26_sva_10_0;
      quad_serial_out_rsci_idat_263 <= for_quad_to_sram_w_z_23_12_sva_11;
      quad_serial_out_rsci_idat_262_252 <= for_quad_to_sram_w_z_23_12_sva_10_0;
      quad_serial_out_rsci_idat_264 <= inputChannel_tmp_7_sva_0;
      quad_serial_out_rsci_idat_276 <= for_inputChannel_tmp_29_sva_11;
      quad_serial_out_rsci_idat_275_265 <= for_inputChannel_tmp_29_sva_10_0;
      quad_serial_out_rsci_idat_288 <= for_quad_to_sram_d_plane_23_12_sva_11;
      quad_serial_out_rsci_idat_287_277 <= for_quad_to_sram_d_plane_23_12_sva_10_0;
      quad_serial_out_rsci_idat_295_289 <= inputChannel_tmp_11_sva_6_0;
      quad_serial_out_rsci_idat_307 <= for_inputChannel_tmp_32_sva_11;
      quad_serial_out_rsci_idat_306_296 <= for_inputChannel_tmp_32_sva_10_0;
      quad_serial_out_rsci_idat_319_308 <= for_quad_to_sram_quad_color_r_23_12_sva;
      quad_serial_out_rsci_idat_322_320 <= for_for_slc_for_inputChannel_tmp_34_2_0_1_itm;
      quad_serial_out_rsci_idat_334 <= for_inputChannel_tmp_35_sva_11;
      quad_serial_out_rsci_idat_333_323 <= for_inputChannel_tmp_35_sva_10_0;
      quad_serial_out_rsci_idat_346_335 <= for_quad_to_sram_quad_color_g_23_12_sva;
      quad_serial_out_rsci_idat_349_347 <= for_for_slc_for_inputChannel_tmp_37_2_0_1_itm;
      quad_serial_out_rsci_idat_361 <= for_inputChannel_tmp_38_sva_11;
      quad_serial_out_rsci_idat_360_350 <= for_inputChannel_tmp_38_sva_10_0;
      quad_serial_out_rsci_idat_373_362 <= for_quad_to_sram_quad_color_b_23_12_sva;
      quad_serial_out_rsci_idat_376_374 <= inputChannel_rsci_idat_mxwt[2:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_accum_params_rsci_idat_10_0_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_12_11_cse <= 2'b00;
      reg_accum_params_rsci_idat_24_13_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_36_25_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_39_37_cse_2_1 <= 2'b00;
      reg_accum_params_rsci_idat_39_37_cse_0 <= 1'b0;
      reg_accum_params_rsci_idat_51_40_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_63_52_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_66_64_cse_2_1 <= 2'b00;
      reg_accum_params_rsci_idat_66_64_cse_0 <= 1'b0;
      reg_accum_params_rsci_idat_78_67_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_90_79_cse <= 12'b000000000000;
      reg_accum_params_rsci_idat_93_91_cse <= 3'b000;
      reg_accum_params_rsci_idat_104_94_cse_10_7 <= 4'b0000;
      reg_accum_params_rsci_idat_104_94_cse_6_0 <= 7'b0000000;
      reg_accum_params_rsci_idat_115_105_cse_10_6 <= 5'b00000;
      reg_accum_params_rsci_idat_115_105_cse_5_0 <= 6'b000000;
      reg_accum_params_rsci_idat_126_116_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_137_127_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_148_138_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_159_149_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_170_160_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_181_171_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_192_182_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_203_193_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_214_204_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_225_215_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_236_226_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_247_237_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_258_248_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_269_259_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_280_270_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_291_281_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_294_292_cse <= 3'b000;
      reg_accum_params_rsci_idat_305_295_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_316_306_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_319_317_cse <= 3'b000;
      reg_accum_params_rsci_idat_330_320_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_341_331_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_344_342_cse_2 <= 1'b0;
      reg_accum_params_rsci_idat_344_342_cse_1_0 <= 2'b00;
      reg_accum_params_rsci_idat_355_345_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_366_356_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_369_367_cse_2 <= 1'b0;
      reg_accum_params_rsci_idat_369_367_cse_1_0 <= 2'b00;
      reg_accum_params_rsci_idat_380_370_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_391_381_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_394_392_cse_2_1 <= 2'b00;
      reg_accum_params_rsci_idat_394_392_cse_0 <= 1'b0;
      reg_accum_params_rsci_idat_405_395_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_416_406_cse <= 11'b00000000000;
      reg_accum_params_rsci_idat_419_417_cse <= 3'b000;
    end
    else if ( accum_params_and_cse ) begin
      reg_accum_params_rsci_idat_10_0_cse <= inputChannel_tmp_sva_10_0;
      reg_accum_params_rsci_idat_12_11_cse <= for_for_slc_for_inputChannel_tmp_13_1_0_1_itm;
      reg_accum_params_rsci_idat_24_13_cse <= for_quad_to_sram_quad_color_r_23_12_sva;
      reg_accum_params_rsci_idat_36_25_cse <= for_inputChannel_tmp_17_sva;
      reg_accum_params_rsci_idat_39_37_cse_2_1 <= inputChannel_tmp_4_sva_2_1;
      reg_accum_params_rsci_idat_39_37_cse_0 <= inputChannel_tmp_4_sva_0;
      reg_accum_params_rsci_idat_51_40_cse <= for_quad_to_sram_quad_color_g_23_12_sva;
      reg_accum_params_rsci_idat_63_52_cse <= for_inputChannel_tmp_14_sva;
      reg_accum_params_rsci_idat_66_64_cse_2_1 <= inputChannel_tmp_7_sva_2_1;
      reg_accum_params_rsci_idat_66_64_cse_0 <= inputChannel_tmp_7_sva_0;
      reg_accum_params_rsci_idat_78_67_cse <= for_quad_to_sram_quad_color_b_23_12_sva;
      reg_accum_params_rsci_idat_90_79_cse <= for_inputChannel_tmp_11_sva;
      reg_accum_params_rsci_idat_93_91_cse <= for_for_slc_for_inputChannel_tmp_34_2_0_1_itm;
      reg_accum_params_rsci_idat_104_94_cse_10_7 <= inputChannel_tmp_11_sva_10_7;
      reg_accum_params_rsci_idat_104_94_cse_6_0 <= inputChannel_tmp_11_sva_6_0;
      reg_accum_params_rsci_idat_115_105_cse_10_6 <= inputChannel_tmp_12_sva_10_6;
      reg_accum_params_rsci_idat_115_105_cse_5_0 <= inputChannel_tmp_12_sva_5_0;
      reg_accum_params_rsci_idat_126_116_cse <= for_inputChannel_tmp_20_sva_10_0;
      reg_accum_params_rsci_idat_137_127_cse <= for_inputChannel_tmp_23_sva_10_0;
      reg_accum_params_rsci_idat_148_138_cse <= for_inputChannel_tmp_26_sva_10_0;
      reg_accum_params_rsci_idat_159_149_cse <= for_inputChannel_tmp_29_sva_10_0;
      reg_accum_params_rsci_idat_170_160_cse <= for_inputChannel_tmp_32_sva_10_0;
      reg_accum_params_rsci_idat_181_171_cse <= for_inputChannel_tmp_35_sva_10_0;
      reg_accum_params_rsci_idat_192_182_cse <= for_inputChannel_tmp_38_sva_10_0;
      reg_accum_params_rsci_idat_203_193_cse <= for_quad_to_sram_corner_pt_x_sva_10_0;
      reg_accum_params_rsci_idat_214_204_cse <= for_quad_to_sram_corner_pt_y_sva_10_0;
      reg_accum_params_rsci_idat_225_215_cse <= for_quad_to_sram_corner_pt_z_sva_10_0;
      reg_accum_params_rsci_idat_236_226_cse <= for_quad_to_sram_d_plane_23_12_sva_10_0;
      reg_accum_params_rsci_idat_247_237_cse <= for_quad_to_sram_normal_x_23_12_sva_10_0;
      reg_accum_params_rsci_idat_258_248_cse <= for_quad_to_sram_normal_y_23_12_sva_10_0;
      reg_accum_params_rsci_idat_269_259_cse <= for_quad_to_sram_normal_z_23_12_sva_10_0;
      reg_accum_params_rsci_idat_280_270_cse <= for_quad_to_sram_u_x_sva_10_0;
      reg_accum_params_rsci_idat_291_281_cse <= for_quad_to_sram_u_y_sva_10_0;
      reg_accum_params_rsci_idat_294_292_cse <= for_for_slc_for_inputChannel_tmp_37_2_0_1_itm;
      reg_accum_params_rsci_idat_305_295_cse <= for_quad_to_sram_u_z_sva_10_0;
      reg_accum_params_rsci_idat_316_306_cse <= for_quad_to_sram_v_x_sva_10_0;
      reg_accum_params_rsci_idat_319_317_cse <= for_for_slc_for_inputChannel_tmp_9_2_0_1_itm;
      reg_accum_params_rsci_idat_330_320_cse <= for_quad_to_sram_v_y_sva_10_0;
      reg_accum_params_rsci_idat_341_331_cse <= for_quad_to_sram_v_z_sva_10_0;
      reg_accum_params_rsci_idat_344_342_cse_2 <= inputChannel_tmp_35_sva_2;
      reg_accum_params_rsci_idat_344_342_cse_1_0 <= inputChannel_tmp_35_sva_1_0;
      reg_accum_params_rsci_idat_355_345_cse <= for_quad_to_sram_w_x_23_12_sva_10_0;
      reg_accum_params_rsci_idat_366_356_cse <= for_quad_to_sram_w_y_23_12_sva_10_0;
      reg_accum_params_rsci_idat_369_367_cse_2 <= inputChannel_tmp_38_sva_2;
      reg_accum_params_rsci_idat_369_367_cse_1_0 <= inputChannel_tmp_38_sva_1_0;
      reg_accum_params_rsci_idat_380_370_cse <= for_quad_to_sram_w_z_23_12_sva_10_0;
      reg_accum_params_rsci_idat_391_381_cse <= inputChannel_tmp_40_sva_10_0;
      reg_accum_params_rsci_idat_394_392_cse_2_1 <= inputChannel_tmp_41_sva_2_1;
      reg_accum_params_rsci_idat_394_392_cse_0 <= inputChannel_tmp_41_sva_0;
      reg_accum_params_rsci_idat_405_395_cse <= inputChannel_tmp_42_sva_10_0;
      reg_accum_params_rsci_idat_416_406_cse <= inputChannel_tmp_43_sva_10_0;
      reg_accum_params_rsci_idat_419_417_cse <= inputChannel_rsci_idat_mxwt[2:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      qbuffer_params_rsci_idat_10_0 <= 11'b00000000000;
      qbuffer_params_rsci_idat_12_11 <= 2'b00;
      qbuffer_params_rsci_idat_23_20 <= 4'b0000;
      qbuffer_params_rsci_idat_19_13 <= 7'b0000000;
      qbuffer_params_rsci_idat_34_30 <= 5'b00000;
      qbuffer_params_rsci_idat_29_24 <= 6'b000000;
      qbuffer_params_rsci_idat_45_35 <= 11'b00000000000;
      qbuffer_params_rsci_idat_56_46 <= 11'b00000000000;
    end
    else if ( qbuffer_params_and_cse ) begin
      qbuffer_params_rsci_idat_10_0 <= inputChannel_tmp_sva_10_0;
      qbuffer_params_rsci_idat_12_11 <= for_for_slc_for_inputChannel_tmp_13_1_0_1_itm;
      qbuffer_params_rsci_idat_23_20 <= inputChannel_tmp_11_sva_10_7;
      qbuffer_params_rsci_idat_19_13 <= inputChannel_tmp_11_sva_6_0;
      qbuffer_params_rsci_idat_34_30 <= inputChannel_tmp_12_sva_10_6;
      qbuffer_params_rsci_idat_29_24 <= inputChannel_tmp_12_sva_5_0;
      qbuffer_params_rsci_idat_45_35 <= for_inputChannel_tmp_20_sva_10_0;
      qbuffer_params_rsci_idat_56_46 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_quad_serial_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_accum_params_rsci_ivld_run_psct_cse <= 1'b0;
      reg_qbuffer_params_rsci_ivld_run_psct_cse <= 1'b0;
      reg_inputChannel_rsci_irdy_run_psct_cse <= 1'b0;
      inputChannel_tmp_43_sva_10_0 <= 11'b00000000000;
    end
    else if ( run_wen ) begin
      reg_quad_serial_out_rsci_ivld_run_psct_cse <= (fsm_output[1]) & (~ (fsm_output[3]))
          & and_380_cse & (fsm_output[6:4]==3'b101);
      reg_accum_params_rsci_ivld_run_psct_cse <= (~ (fsm_output[1])) & (fsm_output[3])
          & and_380_cse & (fsm_output[6:4]==3'b010);
      reg_qbuffer_params_rsci_ivld_run_psct_cse <= and_356_cse & and_380_cse & nor_173_cse
          & (~ (fsm_output[6]));
      reg_inputChannel_rsci_irdy_run_psct_cse <= ~ (mux_117_nl);
      inputChannel_tmp_43_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_sva_10_0 <= 11'b00000000000;
    end
    else if ( run_wen & (mux_120_nl) ) begin
      inputChannel_tmp_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_slc_for_inputChannel_tmp_13_1_0_1_itm <= 2'b00;
    end
    else if ( run_wen & (~((mux_121_nl) | (fsm_output[0]) | (fsm_output[6]))) ) begin
      for_for_slc_for_inputChannel_tmp_13_1_0_1_itm <= inputChannel_rsci_idat_mxwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_quad_color_r_23_12_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~((mux_122_nl) | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[5])))
        ) begin
      for_quad_to_sram_quad_color_r_23_12_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_17_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~(or_314_cse | (fsm_output[0]) | (fsm_output[5]) | (~((fsm_output[2])
        ^ (fsm_output[6]))) | (fsm_output[4]))) ) begin
      for_inputChannel_tmp_17_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_4_sva_2_1 <= 2'b00;
    end
    else if ( (~ (mux_237_nl)) & (~ (fsm_output[5])) & run_wen ) begin
      inputChannel_tmp_4_sva_2_1 <= inputChannel_rsci_idat_mxwt[2:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_4_sva_0 <= 1'b0;
    end
    else if ( (~ (fsm_output[5])) & (fsm_output[2]) & (fsm_output[0]) & (~ (fsm_output[4]))
        & nor_177_cse & run_wen ) begin
      inputChannel_tmp_4_sva_0 <= MUX_s_1_2_2((inputChannel_rsci_idat_mxwt[0]), (inputChannel_rsci_idat_mxwt[0]),
          and_27_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_quad_color_g_23_12_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~((mux_127_nl) | or_dcpl_30)) ) begin
      for_quad_to_sram_quad_color_g_23_12_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_14_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~((mux_128_nl) | nand_44_cse | (fsm_output[6]))) ) begin
      for_inputChannel_tmp_14_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_7_sva_2_1 <= 2'b00;
    end
    else if ( (~ (mux_241_nl)) & (~ (fsm_output[5])) & run_wen ) begin
      inputChannel_tmp_7_sva_2_1 <= inputChannel_rsci_idat_mxwt[2:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_7_sva_0 <= 1'b0;
    end
    else if ( (~((mux_242_nl) | (fsm_output[5]))) & (fsm_output[4:2]==3'b010) & run_wen
        ) begin
      inputChannel_tmp_7_sva_0 <= MUX_s_1_2_2((inputChannel_rsci_idat_mxwt[0]), (inputChannel_rsci_idat_mxwt[0]),
          and_31_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_quad_color_b_23_12_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~((mux_132_nl) | (fsm_output[5]))) ) begin
      for_quad_to_sram_quad_color_b_23_12_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_11_sva <= 12'b000000000000;
    end
    else if ( run_wen & (~(nand_33_cse | (fsm_output[0]) | (fsm_output[2]) | ((fsm_output[5])
        ^ (fsm_output[4])) | (fsm_output[6]))) ) begin
      for_inputChannel_tmp_11_sva <= inputChannel_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_slc_for_inputChannel_tmp_34_2_0_1_itm <= 3'b000;
    end
    else if ( run_wen & (~((mux_133_nl) | or_dcpl_40 | (fsm_output[5]))) ) begin
      for_for_slc_for_inputChannel_tmp_34_2_0_1_itm <= inputChannel_rsci_idat_mxwt[2:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_11_sva_10_7 <= 4'b0000;
    end
    else if ( (mux_244_nl) & (~ (fsm_output[5])) & run_wen ) begin
      inputChannel_tmp_11_sva_10_7 <= inputChannel_rsci_idat_mxwt[10:7];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_11_sva_6_0 <= 7'b0000000;
    end
    else if ( nor_173_cse & (~((fsm_output[1]) ^ (fsm_output[6]))) & (fsm_output[2])
        & (~ (fsm_output[0])) & (fsm_output[3]) & run_wen ) begin
      inputChannel_tmp_11_sva_6_0 <= inputChannel_rsci_idat_mxwt[6:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_12_sva_10_6 <= 5'b00000;
    end
    else if ( (mux_252_nl) & run_wen ) begin
      inputChannel_tmp_12_sva_10_6 <= mux_225_rgt[10:6];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_12_sva_5_0 <= 6'b000000;
    end
    else if ( (mux_253_nl) & (~ (fsm_output[4])) & (fsm_output[2]) & (fsm_output[3])
        & (~ (fsm_output[6])) & run_wen ) begin
      inputChannel_tmp_12_sva_5_0 <= mux_225_rgt[5:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_20_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_257_nl)) & run_wen ) begin
      for_inputChannel_tmp_20_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_20_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_258_nl) & (fsm_output[1]) & (~ (fsm_output[5])) & (~ (fsm_output[4]))
        & run_wen ) begin
      for_inputChannel_tmp_20_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_23_sva_11 <= 1'b0;
    end
    else if ( (mux_260_nl) & run_wen ) begin
      for_inputChannel_tmp_23_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_23_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_261_nl) & (fsm_output[2]) & (fsm_output[1]) & (~ (fsm_output[4]))
        & (~ (fsm_output[5])) & run_wen ) begin
      for_inputChannel_tmp_23_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_26_sva_11 <= 1'b0;
    end
    else if ( (mux_263_nl) & run_wen ) begin
      for_inputChannel_tmp_26_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_26_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_264_nl) & nor_164_cse & (~ (fsm_output[5])) & run_wen ) begin
      for_inputChannel_tmp_26_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_29_sva_11 <= 1'b0;
    end
    else if ( (mux_266_nl) & run_wen ) begin
      for_inputChannel_tmp_29_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_29_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_267_nl) & (~((fsm_output[1]) | (fsm_output[5]))) & run_wen ) begin
      for_inputChannel_tmp_29_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_32_sva_11 <= 1'b0;
    end
    else if ( (mux_269_nl) & run_wen ) begin
      for_inputChannel_tmp_32_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_32_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_270_nl) & (fsm_output[1]) & (~ (fsm_output[5])) & run_wen ) begin
      for_inputChannel_tmp_32_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_35_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_275_nl)) & run_wen ) begin
      for_inputChannel_tmp_35_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_35_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[5:4]==2'b01) & ((fsm_output[0]) ^ (fsm_output[6])) & (fsm_output[3:1]==3'b001)
        & run_wen ) begin
      for_inputChannel_tmp_35_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_38_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_280_nl)) & run_wen ) begin
      for_inputChannel_tmp_38_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_inputChannel_tmp_38_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[5:4]==2'b01) & (~((fsm_output[0]) ^ (fsm_output[6]))) &
        nor_177_cse & (fsm_output[2]) & run_wen ) begin
      for_inputChannel_tmp_38_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_x_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_286_nl)) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_corner_pt_x_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_x_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_287_nl) & (~ (fsm_output[6])) & (fsm_output[2]) & (fsm_output[0])
        & run_wen ) begin
      for_quad_to_sram_corner_pt_x_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_y_sva_11 <= 1'b0;
    end
    else if ( (mux_289_nl) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_corner_pt_y_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_y_sva_10_0 <= 11'b00000000000;
    end
    else if ( mux_290_cse & (fsm_output[4]) & nor_148_cse & (~ (fsm_output[0])) &
        run_wen ) begin
      for_quad_to_sram_corner_pt_y_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_z_sva_11 <= 1'b0;
    end
    else if ( (mux_292_nl) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_corner_pt_z_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_corner_pt_z_sva_10_0 <= 11'b00000000000;
    end
    else if ( mux_290_cse & (fsm_output[4]) & nor_148_cse & (fsm_output[0]) & run_wen
        ) begin
      for_quad_to_sram_corner_pt_z_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_d_plane_23_12_sva_11 <= 1'b0;
    end
    else if ( (mux_295_nl) & run_wen ) begin
      for_quad_to_sram_d_plane_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_d_plane_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_296_nl) & (fsm_output[3]) & (~ (fsm_output[1])) & (~ (fsm_output[5]))
        & run_wen ) begin
      for_quad_to_sram_d_plane_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_x_23_12_sva_11 <= 1'b0;
    end
    else if ( (mux_298_nl) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_normal_x_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_x_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[4]) & (~ (fsm_output[6])) & (~((fsm_output[1]) ^ (fsm_output[5])))
        & (fsm_output[3]) & (fsm_output[0]) & (~ (fsm_output[2])) & run_wen ) begin
      for_quad_to_sram_normal_x_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_y_23_12_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_302_nl)) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_normal_y_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_y_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[4]) & (~ (fsm_output[6])) & (~((fsm_output[2]) ^ (fsm_output[5])))
        & (fsm_output[3]) & (fsm_output[1]) & (~ (fsm_output[0])) & run_wen ) begin
      for_quad_to_sram_normal_y_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_z_23_12_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_306_nl)) & run_wen ) begin
      for_quad_to_sram_normal_z_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_normal_z_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_307_nl) & (fsm_output[0]) & (~ (fsm_output[2])) & (~ (fsm_output[5]))
        & run_wen ) begin
      for_quad_to_sram_normal_z_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_x_sva_11 <= 1'b0;
    end
    else if ( (mux_309_nl) & run_wen & (~ (fsm_output[6])) ) begin
      for_quad_to_sram_u_x_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_x_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_310_nl) & (~ (fsm_output[0])) & (fsm_output[4]) & run_wen & (~
        (fsm_output[6])) ) begin
      for_quad_to_sram_u_x_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_y_sva_11 <= 1'b0;
    end
    else if ( (mux_312_nl) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_u_y_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_y_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_313_nl) & (~ (fsm_output[6])) & (fsm_output[4]) & (fsm_output[0])
        & run_wen ) begin
      for_quad_to_sram_u_y_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_slc_for_inputChannel_tmp_37_2_0_1_itm <= 3'b000;
    end
    else if ( run_wen & (~((fsm_output[0]) | (~ (fsm_output[2])) | or_214_cse | (mux_185_nl)))
        ) begin
      for_for_slc_for_inputChannel_tmp_37_2_0_1_itm <= inputChannel_rsci_idat_mxwt[2:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_z_sva_11 <= 1'b0;
    end
    else if ( (mux_315_nl) & (~ (fsm_output[6])) & run_wen ) begin
      for_quad_to_sram_u_z_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_u_z_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_316_nl) & (fsm_output[2]) & (~ (fsm_output[6])) & run_wen & (fsm_output[4])
        ) begin
      for_quad_to_sram_u_z_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_x_sva_11 <= 1'b0;
    end
    else if ( (mux_317_nl) & (fsm_output[6:5]==2'b01) & run_wen ) begin
      for_quad_to_sram_v_x_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_x_sva_10_0 <= 11'b00000000000;
    end
    else if ( (mux_318_nl) & (fsm_output[5]) & nor_148_cse & (~ (fsm_output[1]))
        & run_wen ) begin
      for_quad_to_sram_v_x_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_slc_for_inputChannel_tmp_9_2_0_1_itm <= 3'b000;
    end
    else if ( run_wen & (~((mux_191_nl) | (fsm_output[1]) | (fsm_output[2]) | (~
        (fsm_output[5])) | (fsm_output[6]))) ) begin
      for_for_slc_for_inputChannel_tmp_9_2_0_1_itm <= inputChannel_rsci_idat_mxwt[2:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_y_sva_11 <= 1'b0;
    end
    else if ( (mux_320_nl) & (fsm_output[6:5]==2'b01) & run_wen ) begin
      for_quad_to_sram_v_y_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_y_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[6:5]==2'b01) & xnor_2_cse & (~ (fsm_output[3])) & (fsm_output[1])
        & (~ (fsm_output[0])) & run_wen ) begin
      for_quad_to_sram_v_y_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_z_sva_11 <= 1'b0;
    end
    else if ( (mux_324_nl) & (fsm_output[6:5]==2'b01) & run_wen ) begin
      for_quad_to_sram_v_z_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_v_z_sva_10_0 <= 11'b00000000000;
    end
    else if ( (fsm_output[6:5]==2'b01) & xnor_2_cse & (~ (fsm_output[3])) & (fsm_output[1])
        & (fsm_output[0]) & run_wen ) begin
      for_quad_to_sram_v_z_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_35_sva_2 <= 1'b0;
    end
    else if ( (mux_326_nl) & run_wen ) begin
      inputChannel_tmp_35_sva_2 <= inputChannel_rsci_idat_mxwt[2];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_35_sva_1_0 <= 2'b00;
    end
    else if ( (mux_327_nl) & (fsm_output[2]) & (~ (fsm_output[6])) & run_wen & (fsm_output[5])
        ) begin
      inputChannel_tmp_35_sva_1_0 <= inputChannel_rsci_idat_mxwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_x_23_12_sva_11 <= 1'b0;
    end
    else if ( (~ (mux_330_nl)) & (~ (fsm_output[4])) & run_wen ) begin
      for_quad_to_sram_w_x_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_x_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (~((mux_331_nl) | (fsm_output[4]))) & (fsm_output[3:1]==3'b010) & run_wen
        ) begin
      for_quad_to_sram_w_x_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_y_23_12_sva_11 <= 1'b0;
    end
    else if ( (mux_335_nl) & (~ (fsm_output[4])) & run_wen ) begin
      for_quad_to_sram_w_y_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_y_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (~((mux_336_nl) | (fsm_output[4]))) & (fsm_output[3:1]==3'b011) & run_wen
        ) begin
      for_quad_to_sram_w_y_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_38_sva_2 <= 1'b0;
    end
    else if ( (mux_339_nl) & run_wen ) begin
      inputChannel_tmp_38_sva_2 <= inputChannel_rsci_idat_mxwt[2];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_38_sva_1_0 <= 2'b00;
    end
    else if ( (mux_340_nl) & (~ (fsm_output[4])) & (fsm_output[1]) & (~ (fsm_output[3]))
        & run_wen ) begin
      inputChannel_tmp_38_sva_1_0 <= inputChannel_rsci_idat_mxwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_z_23_12_sva_11 <= 1'b0;
    end
    else if ( (mux_341_nl) & (fsm_output[4:3]==2'b01) & run_wen ) begin
      for_quad_to_sram_w_z_23_12_sva_11 <= inputChannel_rsci_idat_mxwt[11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_quad_to_sram_w_z_23_12_sva_10_0 <= 11'b00000000000;
    end
    else if ( (~((mux_342_nl) | (fsm_output[4]))) & (fsm_output[3]) & (~ (fsm_output[2]))
        & (~ (fsm_output[0])) & run_wen ) begin
      for_quad_to_sram_w_z_23_12_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_40_sva_10_0 <= 11'b00000000000;
    end
    else if ( run_wen & (~(or_dcpl_69 | or_dcpl_11)) ) begin
      inputChannel_tmp_40_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_41_sva_2_1 <= 2'b00;
    end
    else if ( (mux_344_nl) & run_wen ) begin
      inputChannel_tmp_41_sva_2_1 <= inputChannel_rsci_idat_mxwt[2:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_41_sva_0 <= 1'b0;
    end
    else if ( (~((mux_345_nl) | (fsm_output[4]))) & nor_125_cse & (fsm_output[3])
        & run_wen ) begin
      inputChannel_tmp_41_sva_0 <= MUX_s_1_2_2((inputChannel_rsci_idat_mxwt[0]),
          (inputChannel_rsci_idat_mxwt[0]), and_111_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      inputChannel_tmp_42_sva_10_0 <= 11'b00000000000;
    end
    else if ( run_wen & (~((fsm_output[2]) | (~ and_348_cse) | or_dcpl_11)) ) begin
      inputChannel_tmp_42_sva_10_0 <= inputChannel_rsci_idat_mxwt[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_33_true_operator_33_true_and_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_18 | or_dcpl_11)) ) begin
      operator_33_true_operator_33_true_and_itm <= (inputChannel_tmp_12_sva_5_0 ==
          (operator_11_false_acc_sdt_sva_1[5:0])) & (operator_11_false_acc_sdt_sva_1[11:6]==6'b000000);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_slc_for_acc_6_itm <= 1'b0;
    end
    else if ( run_wen & (mux_219_nl) ) begin
      for_slc_for_acc_6_itm <= readslicef_7_1_6((for_acc_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_slc_for_inputChannel_tmp_10_0_1_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_69 | (~ and_dcpl_61) | (fsm_output[6]))) ) begin
      for_for_slc_for_inputChannel_tmp_10_0_1_itm <= inputChannel_rsci_idat_mxwt[0];
    end
  end
  assign nor_14_nl = ~((fsm_output[5:0]!=6'b101101));
  assign mux_114_nl = MUX_s_1_2_2(and_356_cse, (fsm_output[3]), fsm_output[0]);
  assign mux_113_nl = MUX_s_1_2_2((fsm_output[3]), or_314_cse, fsm_output[0]);
  assign mux_115_nl = MUX_s_1_2_2((mux_114_nl), (mux_113_nl), fsm_output[2]);
  assign or_23_nl = (fsm_output[5]) | (mux_115_nl);
  assign mux_116_nl = MUX_s_1_2_2((fsm_output[5]), (or_23_nl), fsm_output[4]);
  assign mux_117_nl = MUX_s_1_2_2((nor_14_nl), (mux_116_nl), fsm_output[6]);
  assign nor_16_nl = ~((fsm_output[5:1]!=5'b00000));
  assign mux_120_nl = MUX_s_1_2_2((nor_16_nl), mux_tmp_7, fsm_output[6]);
  assign or_31_nl = (fsm_output[5]) | (fsm_output[2]) | (fsm_output[3]) | (~ (fsm_output[1]));
  assign nand_5_nl = ~((fsm_output[5]) & (fsm_output[2]) & (fsm_output[3]) & (~ (fsm_output[1])));
  assign mux_121_nl = MUX_s_1_2_2((or_31_nl), (nand_5_nl), fsm_output[4]);
  assign or_36_nl = (fsm_output[4]) | (~((fsm_output[1:0]==2'b11)));
  assign or_35_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[1]);
  assign mux_122_nl = MUX_s_1_2_2((or_36_nl), (or_35_nl), fsm_output[6]);
  assign or_169_nl = (fsm_output[1]) | (fsm_output[3]) | (fsm_output[4]) | (~ and_380_cse);
  assign nor_178_nl = ~((fsm_output[4]) | and_380_cse);
  assign mux_235_nl = MUX_s_1_2_2((nor_178_nl), (fsm_output[4]), fsm_output[3]);
  assign mux_233_nl = MUX_s_1_2_2((~ (fsm_output[2])), and_380_cse, fsm_output[4]);
  assign mux_234_nl = MUX_s_1_2_2((mux_233_nl), (fsm_output[4]), fsm_output[3]);
  assign mux_236_nl = MUX_s_1_2_2((mux_235_nl), (mux_234_nl), fsm_output[1]);
  assign mux_237_nl = MUX_s_1_2_2((or_169_nl), (mux_236_nl), fsm_output[6]);
  assign mux_124_nl = MUX_s_1_2_2((fsm_output[3]), or_42_cse, fsm_output[2]);
  assign mux_125_nl = MUX_s_1_2_2((mux_124_nl), (~ mux_tmp_11), fsm_output[4]);
  assign and_27_nl = (mux_125_nl) & and_dcpl_26;
  assign or_48_nl = (fsm_output[4]) | (~ (fsm_output[2])) | (fsm_output[0]);
  assign or_47_nl = (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[0]));
  assign mux_127_nl = MUX_s_1_2_2((or_48_nl), (or_47_nl), fsm_output[6]);
  assign or_51_nl = (~ (fsm_output[5])) | (~ (fsm_output[3])) | (fsm_output[1]);
  assign mux_128_nl = MUX_s_1_2_2(or_dcpl_30, (or_51_nl), fsm_output[4]);
  assign or_173_nl = (fsm_output[0]) | (fsm_output[6]) | (fsm_output[4]);
  assign or_172_nl = (~ (fsm_output[0])) | (~ (fsm_output[6])) | (fsm_output[4]);
  assign mux_239_nl = MUX_s_1_2_2((or_173_nl), (or_172_nl), fsm_output[1]);
  assign mux_240_nl = MUX_s_1_2_2(not_tmp_90, (mux_239_nl), fsm_output[3]);
  assign or_171_nl = and_383_cse | not_tmp_90;
  assign or_170_nl = (~ (fsm_output[6])) | (fsm_output[4]);
  assign mux_238_nl = MUX_s_1_2_2((or_171_nl), (or_170_nl), fsm_output[3]);
  assign mux_241_nl = MUX_s_1_2_2((mux_240_nl), (mux_238_nl), fsm_output[2]);
  assign mux_129_nl = MUX_s_1_2_2(and_348_cse, (fsm_output[3]), fsm_output[2]);
  assign mux_130_nl = MUX_s_1_2_2((mux_129_nl), (~ mux_tmp_11), fsm_output[4]);
  assign and_31_nl = (mux_130_nl) & and_dcpl_26;
  assign or_339_nl = (fsm_output[0]) | (fsm_output[6]);
  assign nand_54_nl = ~((fsm_output[0]) & (fsm_output[6]));
  assign mux_242_nl = MUX_s_1_2_2((or_339_nl), (nand_54_nl), fsm_output[1]);
  assign or_57_nl = (fsm_output[4:0]!=5'b01001);
  assign or_56_nl = (fsm_output[4:0]!=5'b10110);
  assign mux_132_nl = MUX_s_1_2_2((or_57_nl), (or_56_nl), fsm_output[6]);
  assign or_66_nl = (fsm_output[4]) | nand_33_cse;
  assign or_65_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[1]);
  assign mux_133_nl = MUX_s_1_2_2((or_66_nl), (or_65_nl), fsm_output[6]);
  assign nor_174_nl = ~((fsm_output[4:0]!=5'b01100));
  assign and_382_nl = nand_53_cse & (fsm_output[4]);
  assign nor_175_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[4]));
  assign mux_243_nl = MUX_s_1_2_2((and_382_nl), (nor_175_nl), fsm_output[3]);
  assign mux_244_nl = MUX_s_1_2_2((nor_174_nl), (mux_243_nl), fsm_output[6]);
  assign mux_249_nl = MUX_s_1_2_2(and_dcpl_61, mux_248_cse, and_380_cse);
  assign mux_247_nl = MUX_s_1_2_2(and_dcpl_61, (fsm_output[5]), fsm_output[2]);
  assign mux_250_nl = MUX_s_1_2_2((mux_249_nl), (mux_247_nl), fsm_output[1]);
  assign mux_251_nl = MUX_s_1_2_2(and_dcpl_61, (mux_250_nl), fsm_output[3]);
  assign or_179_nl = (fsm_output[5:4]!=2'b00);
  assign mux_245_nl = MUX_s_1_2_2((fsm_output[5]), (or_179_nl), or_178_cse);
  assign mux_246_nl = MUX_s_1_2_2((fsm_output[5]), (mux_245_nl), fsm_output[3]);
  assign mux_252_nl = MUX_s_1_2_2((mux_251_nl), (~ (mux_246_nl)), fsm_output[6]);
  assign nor_172_nl = ~((~ (fsm_output[0])) | (fsm_output[5]));
  assign mux_253_nl = MUX_s_1_2_2((nor_172_nl), (fsm_output[5]), fsm_output[1]);
  assign and_378_nl = (fsm_output[3:2]==2'b11);
  assign mux_254_nl = MUX_s_1_2_2(and_131_cse, (and_378_nl), fsm_output[0]);
  assign mux_255_nl = MUX_s_1_2_2((~ and_131_cse), (mux_254_nl), fsm_output[5]);
  assign mux_256_nl = MUX_s_1_2_2((mux_255_nl), (fsm_output[5]), fsm_output[4]);
  assign or_182_nl = (fsm_output[5:0]!=6'b000011);
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), (or_182_nl), fsm_output[6]);
  assign nor_170_nl = ~((fsm_output[0]) | nand_52_cse);
  assign nor_171_nl = ~((~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3]));
  assign mux_258_nl = MUX_s_1_2_2((nor_170_nl), (nor_171_nl), fsm_output[6]);
  assign or_337_nl = (fsm_output[4]) | and_377_cse;
  assign mux_259_nl = MUX_s_1_2_2((or_337_nl), nor_168_cse, fsm_output[5]);
  assign nor_169_nl = ~((fsm_output[5:0]!=6'b000110));
  assign mux_260_nl = MUX_s_1_2_2((mux_259_nl), (nor_169_nl), fsm_output[6]);
  assign and_376_nl = (fsm_output[3]) & (fsm_output[0]);
  assign nor_167_nl = ~((fsm_output[3]) | (fsm_output[0]));
  assign mux_261_nl = MUX_s_1_2_2((and_376_nl), (nor_167_nl), fsm_output[6]);
  assign mux_262_nl = MUX_s_1_2_2((fsm_output[4]), nor_168_cse, fsm_output[5]);
  assign nor_166_nl = ~((fsm_output[5:0]!=6'b001001));
  assign mux_263_nl = MUX_s_1_2_2((mux_262_nl), (nor_166_nl), fsm_output[6]);
  assign nor_162_nl = ~((~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[0]));
  assign nor_163_nl = ~((fsm_output[4]) | (~((fsm_output[3]) & (fsm_output[0]))));
  assign mux_264_nl = MUX_s_1_2_2((nor_162_nl), (nor_163_nl), fsm_output[6]);
  assign and_374_nl = (fsm_output[4]) & ((fsm_output[3:0]!=4'b0000));
  assign mux_265_nl = MUX_s_1_2_2((and_374_nl), nor_168_cse, fsm_output[5]);
  assign nor_161_nl = ~((fsm_output[5]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[1])
      | nand_52_cse);
  assign mux_266_nl = MUX_s_1_2_2((mux_265_nl), (nor_161_nl), fsm_output[6]);
  assign nor_157_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[0])) | (fsm_output[3])
      | (fsm_output[2]));
  assign nor_158_nl = ~((fsm_output[4]) | (fsm_output[0]) | nand_52_cse);
  assign mux_267_nl = MUX_s_1_2_2((nor_157_nl), (nor_158_nl), fsm_output[6]);
  assign and_373_nl = (fsm_output[4]) & ((fsm_output[3:1]!=3'b000));
  assign mux_268_nl = MUX_s_1_2_2((and_373_nl), nor_168_cse, fsm_output[5]);
  assign nor_156_nl = ~((fsm_output[5:0]!=6'b001111));
  assign mux_269_nl = MUX_s_1_2_2((mux_268_nl), (nor_156_nl), fsm_output[6]);
  assign nor_153_nl = ~((~ (fsm_output[4])) | (fsm_output[2]) | (fsm_output[0]) |
      (fsm_output[3]));
  assign nor_154_nl = ~((fsm_output[4]) | (~((fsm_output[2]) & (fsm_output[0]) &
      (fsm_output[3]))));
  assign mux_270_nl = MUX_s_1_2_2((nor_153_nl), (nor_154_nl), fsm_output[6]);
  assign or_215_nl = and_383_cse | (fsm_output[3]);
  assign mux_273_nl = MUX_s_1_2_2(or_216_cse, mux_248_cse, or_215_nl);
  assign mux_274_nl = MUX_s_1_2_2((mux_273_nl), mux_272_cse, fsm_output[2]);
  assign or_212_nl = (fsm_output[5:0]!=6'b010010);
  assign mux_275_nl = MUX_s_1_2_2((mux_274_nl), (or_212_nl), fsm_output[6]);
  assign mux_278_nl = MUX_s_1_2_2(or_216_cse, mux_248_cse, fsm_output[3]);
  assign mux_279_nl = MUX_s_1_2_2((mux_278_nl), mux_272_cse, fsm_output[2]);
  assign or_218_nl = (fsm_output[5:0]!=6'b010101);
  assign mux_280_nl = MUX_s_1_2_2((mux_279_nl), (or_218_nl), fsm_output[6]);
  assign and_368_nl = or_338_cse & (fsm_output[2]);
  assign mux_285_nl = MUX_s_1_2_2(or_216_cse, mux_tmp_160, and_368_nl);
  assign mux_283_nl = MUX_s_1_2_2(mux_tmp_160, or_214_cse, and_369_cse);
  assign nor_62_nl = ~((fsm_output[2:1]!=2'b10));
  assign mux_282_nl = MUX_s_1_2_2(mux_tmp_160, or_214_cse, nor_62_nl);
  assign mux_284_nl = MUX_s_1_2_2((mux_283_nl), (mux_282_nl), fsm_output[0]);
  assign mux_286_nl = MUX_s_1_2_2((mux_285_nl), (mux_284_nl), fsm_output[3]);
  assign nor_150_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[5]));
  assign nor_151_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (~ (fsm_output[5])));
  assign mux_287_nl = MUX_s_1_2_2((nor_150_nl), (nor_151_nl), fsm_output[3]);
  assign and_365_nl = (and_369_cse | (fsm_output[3])) & (fsm_output[4]);
  assign nand_46_nl = ~(or_42_cse & (fsm_output[4]));
  assign mux_288_nl = MUX_s_1_2_2((nand_46_nl), nor_149_cse, fsm_output[2]);
  assign mux_289_nl = MUX_s_1_2_2((and_365_nl), (mux_288_nl), fsm_output[5]);
  assign and_361_nl = or_326_cse & (fsm_output[4]);
  assign nand_45_nl = ~(((~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[3]))
      & (fsm_output[4]));
  assign mux_291_nl = MUX_s_1_2_2((nand_45_nl), nor_149_cse, fsm_output[2]);
  assign mux_292_nl = MUX_s_1_2_2((and_361_nl), (mux_291_nl), fsm_output[5]);
  assign and_359_nl = (fsm_output[4:3]==2'b11);
  assign mux_294_nl = MUX_s_1_2_2((and_359_nl), nor_168_cse, fsm_output[5]);
  assign nor_143_nl = ~((fsm_output[5:0]!=6'b001101));
  assign mux_295_nl = MUX_s_1_2_2((mux_294_nl), (nor_143_nl), fsm_output[6]);
  assign nor_140_nl = ~((~ (fsm_output[4])) | (fsm_output[2]) | (fsm_output[0]));
  assign nor_141_nl = ~((fsm_output[4]) | nand_44_cse);
  assign mux_296_nl = MUX_s_1_2_2((nor_140_nl), (nor_141_nl), fsm_output[6]);
  assign and_357_nl = or_178_cse & (fsm_output[4:3]==2'b11);
  assign nand_42_nl = ~((~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[3])))
      & (fsm_output[4]));
  assign mux_297_nl = MUX_s_1_2_2((nand_42_nl), nor_149_cse, fsm_output[2]);
  assign mux_298_nl = MUX_s_1_2_2((and_357_nl), (mux_297_nl), fsm_output[5]);
  assign nand_41_nl = ~(((fsm_output[2:1]!=2'b00)) & (fsm_output[4:3]==2'b11));
  assign mux_299_nl = MUX_s_1_2_2((fsm_output[4]), (~ (fsm_output[4])), and_356_cse);
  assign or_248_nl = (fsm_output[4:3]!=2'b00);
  assign mux_300_nl = MUX_s_1_2_2((mux_299_nl), (or_248_nl), fsm_output[0]);
  assign mux_301_nl = MUX_s_1_2_2((fsm_output[4]), (mux_300_nl), fsm_output[2]);
  assign mux_302_nl = MUX_s_1_2_2((nand_41_nl), (mux_301_nl), fsm_output[5]);
  assign nand_39_nl = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]));
  assign nand_40_nl = ~((fsm_output[4:3]==2'b11));
  assign mux_304_nl = MUX_s_1_2_2((nand_39_nl), (nand_40_nl), fsm_output[2]);
  assign or_252_nl = and_372_cse | (fsm_output[4]);
  assign mux_303_nl = MUX_s_1_2_2((fsm_output[4]), (or_252_nl), fsm_output[2]);
  assign mux_305_nl = MUX_s_1_2_2((mux_304_nl), (mux_303_nl), fsm_output[5]);
  assign or_250_nl = (fsm_output[5:0]!=6'b000001);
  assign mux_306_nl = MUX_s_1_2_2((mux_305_nl), (or_250_nl), fsm_output[6]);
  assign mux_307_nl = MUX_s_1_2_2(and_354_cse, nor_138_cse, fsm_output[6]);
  assign and_353_nl = (fsm_output[4:2]==3'b111);
  assign nor_137_nl = ~((fsm_output[3:0]!=4'b0010));
  assign mux_308_nl = MUX_s_1_2_2(nand_38_cse, (nor_137_nl), fsm_output[4]);
  assign mux_309_nl = MUX_s_1_2_2((and_353_nl), (mux_308_nl), fsm_output[5]);
  assign nor_135_nl = ~((fsm_output[1]) | nand_52_cse);
  assign nor_136_nl = ~((fsm_output[3:1]!=3'b001));
  assign mux_310_nl = MUX_s_1_2_2((nor_135_nl), (nor_136_nl), fsm_output[5]);
  assign and_385_nl = (~(((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[3]))
      & (fsm_output[4]))) & (fsm_output[5]);
  assign nor_133_nl = ~((fsm_output[5:4]!=2'b10));
  assign nor_134_nl = ~((fsm_output[5:4]!=2'b01));
  assign mux_311_nl = MUX_s_1_2_2((nor_133_nl), (nor_134_nl), and_372_cse);
  assign mux_312_nl = MUX_s_1_2_2((and_385_nl), (mux_311_nl), fsm_output[2]);
  assign nor_130_nl = ~((~ (fsm_output[1])) | (fsm_output[3]) | (~ (fsm_output[5])));
  assign nor_131_nl = ~((fsm_output[1]) | (~ (fsm_output[3])) | (fsm_output[5]));
  assign mux_313_nl = MUX_s_1_2_2((nor_130_nl), (nor_131_nl), fsm_output[2]);
  assign mux_185_nl = MUX_s_1_2_2(nand_33_cse, or_314_cse, fsm_output[6]);
  assign and_349_nl = (fsm_output[5]) & nand_38_cse;
  assign nor_129_nl = ~((fsm_output[3:0]!=4'b0100));
  assign mux_314_nl = MUX_s_1_2_2(and_377_cse, (nor_129_nl), fsm_output[5]);
  assign mux_315_nl = MUX_s_1_2_2((and_349_nl), (mux_314_nl), fsm_output[4]);
  assign nor_128_nl = ~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3]));
  assign mux_316_nl = MUX_s_1_2_2(and_348_cse, (nor_128_nl), fsm_output[5]);
  assign nor_127_nl = ~((fsm_output[3:0]!=4'b0101));
  assign mux_317_nl = MUX_s_1_2_2(nand_38_cse, (nor_127_nl), fsm_output[4]);
  assign mux_318_nl = MUX_s_1_2_2(nor_125_cse, and_380_cse, fsm_output[4]);
  assign or_127_nl = (~ (fsm_output[0])) | (fsm_output[3]);
  assign or_126_nl = (fsm_output[0]) | (~ (fsm_output[3]));
  assign mux_191_nl = MUX_s_1_2_2((or_127_nl), (or_126_nl), fsm_output[4]);
  assign nand_34_nl = ~(or_338_cse & (fsm_output[3]));
  assign mux_319_nl = MUX_s_1_2_2(or_314_cse, (nand_34_nl), fsm_output[2]);
  assign nor_124_nl = ~((fsm_output[3:0]!=4'b0110));
  assign mux_320_nl = MUX_s_1_2_2((mux_319_nl), (nor_124_nl), fsm_output[4]);
  assign mux_322_nl = MUX_s_1_2_2((fsm_output[3]), nand_33_cse, fsm_output[2]);
  assign mux_321_nl = MUX_s_1_2_2(nor_177_cse, (fsm_output[3]), fsm_output[2]);
  assign mux_323_nl = MUX_s_1_2_2((mux_322_nl), (~ (mux_321_nl)), fsm_output[0]);
  assign and_346_nl = (fsm_output[3:0]==4'b0111);
  assign mux_324_nl = MUX_s_1_2_2((mux_323_nl), (and_346_nl), fsm_output[4]);
  assign and_344_nl = (fsm_output[6]) & (~(or_326_cse & (fsm_output[4])));
  assign or_313_nl = (fsm_output[4:1]!=4'b0010);
  assign nand_32_nl = ~((fsm_output[4:1]==4'b1111));
  assign mux_325_nl = MUX_s_1_2_2((or_313_nl), (nand_32_nl), fsm_output[0]);
  assign nor_122_nl = ~((fsm_output[6]) | (mux_325_nl));
  assign mux_326_nl = MUX_s_1_2_2((and_344_nl), (nor_122_nl), fsm_output[5]);
  assign mux_327_nl = MUX_s_1_2_2(nor_138_cse, and_354_cse, fsm_output[0]);
  assign mux_329_nl = MUX_s_1_2_2(or_285_cse, or_311_cse, or_338_cse);
  assign nand_24_nl = ~((fsm_output[2]) & (~ (mux_329_nl)));
  assign or_282_nl = (fsm_output[1]) | (fsm_output[0]) | (fsm_output[6]) | (~ (fsm_output[5]));
  assign mux_328_nl = MUX_s_1_2_2(or_311_cse, (or_282_nl), fsm_output[2]);
  assign mux_330_nl = MUX_s_1_2_2((nand_24_nl), (mux_328_nl), fsm_output[3]);
  assign mux_331_nl = MUX_s_1_2_2(or_285_cse, or_311_cse, fsm_output[0]);
  assign mux_332_nl = MUX_s_1_2_2((fsm_output[3]), (~ (fsm_output[3])), fsm_output[1]);
  assign nor_nl = ~((~ (fsm_output[1])) | (fsm_output[3]));
  assign mux_333_nl = MUX_s_1_2_2((mux_332_nl), (nor_nl), fsm_output[0]);
  assign mux_334_nl = MUX_s_1_2_2((fsm_output[3]), (mux_333_nl), fsm_output[2]);
  assign and_342_nl = (fsm_output[5]) & (mux_334_nl);
  assign nor_119_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | (~ (fsm_output[0]))
      | (~ (fsm_output[1])) | (fsm_output[3]));
  assign mux_335_nl = MUX_s_1_2_2((and_342_nl), (nor_119_nl), fsm_output[6]);
  assign or_308_nl = (~ (fsm_output[5])) | (fsm_output[0]);
  assign or_309_nl = (fsm_output[5]) | (~ (fsm_output[0]));
  assign mux_336_nl = MUX_s_1_2_2((or_308_nl), (or_309_nl), fsm_output[6]);
  assign nor_115_nl = ~((fsm_output[5:0]!=6'b100111));
  assign nor_117_nl = ~((fsm_output[2]) | (fsm_output[4]));
  assign and_341_nl = (fsm_output[0]) & (fsm_output[2]) & (fsm_output[4]);
  assign mux_337_nl = MUX_s_1_2_2((nor_117_nl), (and_341_nl), fsm_output[1]);
  assign mux_338_nl = MUX_s_1_2_2((mux_337_nl), (fsm_output[4]), fsm_output[3]);
  assign nor_116_nl = ~((fsm_output[5]) | (mux_338_nl));
  assign mux_339_nl = MUX_s_1_2_2((nor_115_nl), (nor_116_nl), fsm_output[6]);
  assign and_340_nl = (fsm_output[5]) & (fsm_output[0]) & (fsm_output[2]);
  assign nor_114_nl = ~((fsm_output[5]) | (fsm_output[0]) | (fsm_output[2]));
  assign mux_340_nl = MUX_s_1_2_2((and_340_nl), (nor_114_nl), fsm_output[6]);
  assign and_339_nl = (fsm_output[5]) & (~(or_338_cse & (fsm_output[2])));
  assign nor_113_nl = ~((fsm_output[5]) | (fsm_output[0]) | (~ (fsm_output[1])) |
      (fsm_output[2]));
  assign mux_341_nl = MUX_s_1_2_2((and_339_nl), (nor_113_nl), fsm_output[6]);
  assign or_305_nl = (~ (fsm_output[5])) | (fsm_output[1]);
  assign or_306_nl = (fsm_output[5]) | (~ (fsm_output[1]));
  assign mux_342_nl = MUX_s_1_2_2((or_305_nl), (or_306_nl), fsm_output[6]);
  assign nor_110_nl = ~((fsm_output[5:0]!=6'b101010));
  assign nand_28_nl = ~(nand_53_cse & (fsm_output[4]));
  assign mux_343_nl = MUX_s_1_2_2((nand_28_nl), (fsm_output[4]), fsm_output[3]);
  assign nor_111_nl = ~((fsm_output[5]) | (mux_343_nl));
  assign mux_344_nl = MUX_s_1_2_2((nor_110_nl), (nor_111_nl), fsm_output[6]);
  assign mux_212_nl = MUX_s_1_2_2((fsm_output[3]), (~ mux_tmp_11), fsm_output[4]);
  assign and_111_nl = (mux_212_nl) & and_dcpl_26;
  assign nand_27_nl = ~((fsm_output[5]) & (fsm_output[1]));
  assign or_304_nl = (fsm_output[5]) | (fsm_output[1]);
  assign mux_345_nl = MUX_s_1_2_2((nand_27_nl), (or_304_nl), fsm_output[6]);
  assign nl_for_acc_nl = ({1'b1 , for_i_5_0_sva_1_mx0w1}) + 7'b0000001;
  assign for_acc_nl = nl_for_acc_nl[6:0];
  assign or_155_nl = (fsm_output[5]) | (fsm_output[3]);
  assign mux_218_nl = MUX_s_1_2_2((fsm_output[5]), (or_155_nl), fsm_output[4]);
  assign mux_219_nl = MUX_s_1_2_2((~ and_dcpl_61), (mux_218_nl), fsm_output[6]);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64_run
// ------------------------------------------------------------------


module QuadBuffer_64_run (
  clk, arst_n, quads_in_rsc_dat, quads_in_rsc_vld, quads_in_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, quads_out_rsc_dat, quads_out_rsc_vld, quads_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [376:0] quads_in_rsc_dat;
  input quads_in_rsc_vld;
  output quads_in_rsc_rdy;
  input [56:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [376:0] quads_out_rsc_dat;
  output quads_out_rsc_vld;
  input quads_out_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire quads_in_rsci_wen_comp;
  wire [376:0] quads_in_rsci_idat_mxwt;
  wire paramsIn_rsci_wen_comp;
  wire [45:0] paramsIn_rsci_idat_mxwt;
  wire quads_out_rsci_wen_comp;
  reg [24:0] quads_out_rsci_idat_376_352;
  reg [1:0] quads_out_rsci_idat_351_350;
  reg [26:0] quads_out_rsci_idat_349_323;
  reg [2:0] quads_out_rsci_idat_322_320;
  reg [23:0] quads_out_rsci_idat_319_296;
  reg [7:0] quads_out_rsci_idat_295_288;
  reg [22:0] quads_out_rsci_idat_287_265;
  reg [8:0] quads_out_rsci_idat_264_256;
  reg [15:0] quads_out_rsci_idat_255_240;
  reg [15:0] quads_out_rsci_idat_239_224;
  reg [8:0] quads_out_rsci_idat_223_215;
  reg [22:0] quads_out_rsci_idat_214_192;
  reg [1:0] quads_out_rsci_idat_191_190;
  reg [25:0] quads_out_rsci_idat_189_164;
  reg [3:0] quads_out_rsci_idat_163_160;
  reg [21:0] quads_out_rsci_idat_159_138;
  reg [9:0] quads_out_rsci_idat_137_128;
  reg [15:0] quads_out_rsci_idat_127_112;
  reg quads_out_rsci_idat_111;
  reg [2:0] quads_out_rsci_idat_110_108;
  reg [11:0] quads_out_rsci_idat_107_96;
  reg [11:0] quads_out_rsci_idat_95_84;
  reg [11:0] quads_out_rsci_idat_83_72;
  reg [7:0] quads_out_rsci_idat_71_64;
  reg [3:0] quads_out_rsci_idat_63_60;
  reg [11:0] quads_out_rsci_idat_59_48;
  reg [11:0] quads_out_rsci_idat_47_36;
  reg [3:0] quads_out_rsci_idat_35_32;
  reg [7:0] quads_out_rsci_idat_31_24;
  reg [11:0] quads_out_rsci_idat_23_12;
  reg [11:0] quads_out_rsci_idat_11_0;
  wire [1:0] for_1_for_1_and_4_tmp;
  wire [1:0] for_1_mux1h_2098_tmp;
  wire operator_33_true_operator_33_true_or_tmp;
  wire [6:0] for_acc_1_tmp;
  wire [7:0] nl_for_acc_1_tmp;
  wire operator_33_true_equal_tmp;
  wire operator_33_true_operator_33_true_and_tmp;
  wire for_1_for_1_if_and_tmp;
  wire for_1_for_if_for_1_for_if_or_tmp;
  wire [6:0] operator_7_false_acc_tmp;
  wire [7:0] nl_operator_7_false_acc_tmp;
  wire for_1_for_if_unequal_tmp;
  wire [11:0] operator_11_false_2_acc_tmp;
  wire [12:0] nl_operator_11_false_2_acc_tmp;
  wire for_1_for_for_1_for_and_1_tmp;
  wire for_1_for_for_1_for_and_tmp;
  wire for_1_for_1_and_2_tmp;
  wire for_1_for_1_and_1_tmp;
  wire for_and_59_tmp;
  wire for_and_58_tmp;
  wire for_and_57_tmp;
  wire for_and_56_tmp;
  wire for_and_55_tmp;
  wire for_and_54_tmp;
  wire for_and_53_tmp;
  wire for_and_52_tmp;
  wire for_and_51_tmp;
  wire for_and_50_tmp;
  wire for_and_49_tmp;
  wire for_and_48_tmp;
  wire for_and_47_tmp;
  wire for_and_46_tmp;
  wire for_and_45_tmp;
  wire for_and_44_tmp;
  wire for_and_43_tmp;
  wire for_and_42_tmp;
  wire for_and_41_tmp;
  wire for_and_40_tmp;
  wire for_and_39_tmp;
  wire for_and_38_tmp;
  wire for_and_37_tmp;
  wire for_and_36_tmp;
  wire for_and_35_tmp;
  wire for_and_34_tmp;
  wire for_and_33_tmp;
  wire for_and_32_tmp;
  wire for_and_31_tmp;
  wire for_and_30_tmp;
  wire for_and_29_tmp;
  wire for_and_28_tmp;
  wire for_and_27_tmp;
  wire for_and_26_tmp;
  wire for_and_25_tmp;
  wire for_and_24_tmp;
  wire for_and_23_tmp;
  wire for_and_22_tmp;
  wire for_and_21_tmp;
  wire for_and_20_tmp;
  wire for_and_19_tmp;
  wire for_and_18_tmp;
  wire for_and_17_tmp;
  wire for_and_16_tmp;
  wire for_and_15_tmp;
  wire for_and_14_tmp;
  wire for_and_13_tmp;
  wire for_for_nor_tmp;
  wire for_and_11_tmp;
  wire for_and_10_tmp;
  wire for_and_9_tmp;
  wire for_and_8_tmp;
  wire for_and_7_tmp;
  wire for_and_6_tmp;
  wire for_and_5_tmp;
  wire for_and_4_tmp;
  wire for_and_2_tmp;
  wire for_and_1_tmp;
  wire for_and_tmp;
  wire for_1_for_1_or_tmp;
  wire [5:0] for_1_for_1_mux_76_tmp;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire or_tmp_5;
  wire nor_tmp_2;
  wire mux_tmp_2;
  wire mux_tmp_9;
  wire mux_tmp_10;
  wire mux_tmp_11;
  wire mux_tmp_12;
  wire mux_tmp_13;
  wire mux_tmp_14;
  wire mux_tmp_15;
  wire mux_tmp_16;
  wire mux_tmp_17;
  wire mux_tmp_18;
  wire mux_tmp_19;
  wire mux_tmp_20;
  wire mux_tmp_21;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire mux_tmp_24;
  wire mux_tmp_25;
  wire mux_tmp_26;
  wire mux_tmp_27;
  wire mux_tmp_28;
  wire mux_tmp_29;
  wire mux_tmp_30;
  wire mux_tmp_31;
  wire mux_tmp_32;
  wire mux_tmp_33;
  wire mux_tmp_34;
  wire mux_tmp_35;
  wire mux_tmp_36;
  wire mux_tmp_37;
  wire mux_tmp_38;
  wire mux_tmp_39;
  wire mux_tmp_40;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire mux_tmp_43;
  wire mux_tmp_44;
  wire mux_tmp_45;
  wire mux_tmp_46;
  wire mux_tmp_47;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire mux_tmp_51;
  wire mux_tmp_52;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire mux_tmp_58;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire mux_tmp_65;
  wire mux_tmp_66;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire or_tmp_161;
  wire or_tmp_162;
  wire or_dcpl_2;
  wire or_dcpl_12;
  wire or_dcpl_13;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_18;
  wire or_dcpl_21;
  wire or_dcpl_24;
  wire or_dcpl_27;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_35;
  wire or_dcpl_36;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire or_dcpl_47;
  wire or_dcpl_48;
  wire or_dcpl_53;
  wire or_dcpl_58;
  wire or_dcpl_63;
  wire or_dcpl_68;
  wire or_dcpl_69;
  wire or_dcpl_74;
  wire or_dcpl_79;
  wire or_dcpl_84;
  wire or_dcpl_89;
  wire or_dcpl_90;
  wire or_dcpl_95;
  wire or_dcpl_100;
  wire or_dcpl_105;
  reg reg_quads_out_rsci_oswt_cse;
  wire quads_out_and_cse;
  reg reg_paramsIn_rsci_oswt_cse;
  reg reg_quads_in_rsci_oswt_cse;
  reg for_1_or_tmp_1;
  wire [1:0] paramsIn_crt_lpi_1_dfm_12_0_mx0_12_11;
  reg [42:0] for_1_read_request_lpi_1;
  wire [24:0] tot_samples_in_img_mul_psp_sva_1;
  wire [27:0] nl_tot_samples_in_img_mul_psp_sva_1;
  reg [24:0] tot_samples_in_img_mul_psp_lpi_1;
  reg exitL_exitL_exit_for_1_for_lpi_1;
  reg sfi_exit_for_1_lpi_1;
  reg [5:0] for_i_6_0_lpi_1_dfm_1_5_0;
  reg [1:0] lfst_exit_for_1_lpi_1_dfm_1;
  reg main_stage_0_2;
  reg exitL_exit_for_1_sva;
  reg lfst_exitL_exit_for_1_for_lpi_1;
  reg for_1_asn_sft_lpi_1;
  reg for_1_and_1898_itm_1;
  reg main_stage_0_3;
  wire for_1_asn_sft_lpi_1_dfm_mx0;
  wire mux_89_cse;
  wire or_281_tmp;
  wire [42:0] z_out;
  reg [11:0] buffer_bank0_data_31_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_31_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_31_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_32_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_32_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_32_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_30_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_30_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_30_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_33_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_33_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_33_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_29_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_29_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_29_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_34_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_34_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_34_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_28_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_28_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_28_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_35_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_35_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_35_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_27_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_27_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_27_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_36_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_36_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_36_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_26_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_26_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_26_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_37_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_37_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_37_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_25_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_25_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_25_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_38_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_38_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_38_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_24_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_24_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_24_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_39_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_39_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_39_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_23_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_23_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_23_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_40_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_40_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_40_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_22_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_22_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_22_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_41_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_41_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_41_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_21_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_21_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_21_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_42_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_42_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_42_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_20_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_20_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_20_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_43_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_43_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_43_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_19_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_19_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_19_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_44_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_44_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_44_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_18_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_18_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_18_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_45_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_45_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_45_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_17_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_17_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_17_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_46_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_46_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_46_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_16_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_16_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_16_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_47_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_47_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_47_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_15_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_15_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_15_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_48_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_48_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_48_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_14_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_14_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_14_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_49_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_49_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_49_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_13_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_13_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_13_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_50_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_50_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_50_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_12_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_12_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_12_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_51_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_51_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_51_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_11_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_11_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_11_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_52_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_52_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_52_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_10_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_10_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_10_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_53_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_53_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_53_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_9_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_9_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_9_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_54_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_54_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_54_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_8_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_8_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_8_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_55_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_55_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_55_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_7_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_7_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_7_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_56_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_56_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_56_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_6_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_6_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_6_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_57_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_57_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_57_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_5_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_5_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_5_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_58_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_58_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_58_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_4_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_4_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_4_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_59_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_59_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_59_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_3_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_3_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_3_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_60_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_60_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_60_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_2_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_2_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_2_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_61_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_61_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_61_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_1_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_1_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_1_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_62_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_62_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_62_31_24_lpi_1;
  reg [11:0] buffer_bank0_data_0_23_12_lpi_1;
  reg [11:0] buffer_bank0_data_0_11_0_lpi_1;
  reg [7:0] buffer_bank0_data_0_31_24_lpi_1;
  reg [11:0] buffer_bank1_data_31_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_31_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_31_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_31_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_32_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_32_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_32_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_32_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_30_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_30_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_30_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_30_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_33_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_33_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_33_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_33_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_29_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_29_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_29_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_29_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_34_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_34_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_34_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_34_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_28_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_28_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_28_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_28_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_35_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_35_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_35_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_35_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_27_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_27_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_27_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_27_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_36_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_36_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_36_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_36_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_26_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_26_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_26_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_26_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_37_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_37_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_37_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_37_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_25_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_25_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_25_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_25_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_38_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_38_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_38_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_38_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_24_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_24_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_24_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_24_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_39_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_39_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_39_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_39_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_23_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_23_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_23_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_23_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_40_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_40_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_40_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_40_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_22_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_22_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_22_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_22_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_41_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_41_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_41_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_41_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_21_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_21_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_21_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_21_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_42_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_42_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_42_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_42_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_20_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_20_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_20_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_20_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_43_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_43_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_43_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_43_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_19_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_19_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_19_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_19_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_44_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_44_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_44_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_44_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_18_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_18_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_18_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_18_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_45_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_45_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_45_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_45_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_17_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_17_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_17_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_17_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_46_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_46_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_46_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_46_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_16_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_16_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_16_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_16_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_47_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_47_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_47_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_47_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_15_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_15_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_15_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_15_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_48_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_48_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_48_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_48_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_14_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_14_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_14_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_14_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_49_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_49_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_49_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_49_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_13_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_13_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_13_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_13_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_50_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_50_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_50_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_50_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_12_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_12_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_12_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_12_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_51_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_51_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_51_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_51_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_11_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_11_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_11_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_11_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_52_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_52_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_52_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_52_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_10_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_10_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_10_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_10_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_53_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_53_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_53_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_53_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_9_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_9_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_9_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_9_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_54_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_54_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_54_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_54_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_8_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_8_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_8_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_8_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_55_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_55_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_55_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_55_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_7_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_7_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_7_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_7_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_56_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_56_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_56_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_56_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_6_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_6_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_6_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_6_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_57_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_57_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_57_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_57_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_5_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_5_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_5_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_5_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_58_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_58_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_58_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_58_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_4_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_4_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_4_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_4_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_59_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_59_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_59_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_59_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_3_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_3_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_3_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_3_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_60_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_60_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_60_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_60_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_2_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_2_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_2_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_2_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_61_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_61_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_61_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_61_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_1_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_1_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_1_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_1_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_62_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_62_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_62_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_62_31_28_lpi_1;
  reg [11:0] buffer_bank1_data_0_15_4_lpi_1;
  reg [11:0] buffer_bank1_data_0_27_16_lpi_1;
  reg [3:0] buffer_bank1_data_0_3_0_lpi_1;
  reg [3:0] buffer_bank1_data_0_31_28_lpi_1;
  reg [11:0] buffer_bank2_data_31_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_31_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_31_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_32_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_32_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_32_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_30_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_30_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_30_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_33_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_33_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_33_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_29_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_29_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_29_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_34_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_34_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_34_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_28_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_28_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_28_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_35_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_35_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_35_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_27_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_27_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_27_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_36_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_36_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_36_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_26_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_26_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_26_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_37_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_37_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_37_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_25_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_25_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_25_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_38_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_38_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_38_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_24_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_24_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_24_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_39_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_39_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_39_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_23_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_23_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_23_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_40_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_40_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_40_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_22_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_22_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_22_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_41_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_41_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_41_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_21_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_21_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_21_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_42_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_42_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_42_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_20_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_20_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_20_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_43_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_43_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_43_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_19_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_19_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_19_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_44_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_44_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_44_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_18_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_18_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_18_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_45_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_45_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_45_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_17_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_17_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_17_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_46_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_46_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_46_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_16_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_16_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_16_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_47_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_47_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_47_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_15_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_15_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_15_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_48_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_48_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_48_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_14_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_14_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_14_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_49_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_49_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_49_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_13_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_13_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_13_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_50_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_50_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_50_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_12_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_12_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_12_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_51_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_51_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_51_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_11_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_11_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_11_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_52_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_52_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_52_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_10_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_10_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_10_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_53_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_53_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_53_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_9_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_9_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_9_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_54_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_54_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_54_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_8_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_8_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_8_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_55_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_55_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_55_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_7_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_7_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_7_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_56_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_56_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_56_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_6_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_6_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_6_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_57_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_57_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_57_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_5_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_5_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_5_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_58_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_58_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_58_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_4_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_4_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_4_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_59_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_59_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_59_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_3_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_3_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_3_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_60_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_60_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_60_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_2_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_2_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_2_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_61_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_61_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_61_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_1_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_1_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_1_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_62_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_62_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_62_31_20_lpi_1;
  reg [11:0] buffer_bank2_data_0_19_8_lpi_1;
  reg [7:0] buffer_bank2_data_0_7_0_lpi_1;
  reg [11:0] buffer_bank2_data_0_31_20_lpi_1;
  reg [2:0] buffer_bank3_data_31_14_12_lpi_1;
  reg buffer_bank3_data_31_15_lpi_1;
  reg [11:0] buffer_bank3_data_31_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_31_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_32_14_12_lpi_1;
  reg buffer_bank3_data_32_15_lpi_1;
  reg [11:0] buffer_bank3_data_32_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_32_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_30_14_12_lpi_1;
  reg buffer_bank3_data_30_15_lpi_1;
  reg [11:0] buffer_bank3_data_30_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_30_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_33_14_12_lpi_1;
  reg buffer_bank3_data_33_15_lpi_1;
  reg [11:0] buffer_bank3_data_33_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_33_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_29_14_12_lpi_1;
  reg buffer_bank3_data_29_15_lpi_1;
  reg [11:0] buffer_bank3_data_29_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_29_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_34_14_12_lpi_1;
  reg buffer_bank3_data_34_15_lpi_1;
  reg [11:0] buffer_bank3_data_34_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_34_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_28_14_12_lpi_1;
  reg buffer_bank3_data_28_15_lpi_1;
  reg [11:0] buffer_bank3_data_28_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_28_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_35_14_12_lpi_1;
  reg buffer_bank3_data_35_15_lpi_1;
  reg [11:0] buffer_bank3_data_35_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_35_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_27_14_12_lpi_1;
  reg buffer_bank3_data_27_15_lpi_1;
  reg [11:0] buffer_bank3_data_27_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_27_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_36_14_12_lpi_1;
  reg buffer_bank3_data_36_15_lpi_1;
  reg [11:0] buffer_bank3_data_36_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_36_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_26_14_12_lpi_1;
  reg buffer_bank3_data_26_15_lpi_1;
  reg [11:0] buffer_bank3_data_26_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_26_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_37_14_12_lpi_1;
  reg buffer_bank3_data_37_15_lpi_1;
  reg [11:0] buffer_bank3_data_37_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_37_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_25_14_12_lpi_1;
  reg buffer_bank3_data_25_15_lpi_1;
  reg [11:0] buffer_bank3_data_25_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_25_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_38_14_12_lpi_1;
  reg buffer_bank3_data_38_15_lpi_1;
  reg [11:0] buffer_bank3_data_38_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_38_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_24_14_12_lpi_1;
  reg buffer_bank3_data_24_15_lpi_1;
  reg [11:0] buffer_bank3_data_24_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_24_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_39_14_12_lpi_1;
  reg buffer_bank3_data_39_15_lpi_1;
  reg [11:0] buffer_bank3_data_39_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_39_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_23_14_12_lpi_1;
  reg buffer_bank3_data_23_15_lpi_1;
  reg [11:0] buffer_bank3_data_23_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_23_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_40_14_12_lpi_1;
  reg buffer_bank3_data_40_15_lpi_1;
  reg [11:0] buffer_bank3_data_40_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_40_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_22_14_12_lpi_1;
  reg buffer_bank3_data_22_15_lpi_1;
  reg [11:0] buffer_bank3_data_22_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_22_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_41_14_12_lpi_1;
  reg buffer_bank3_data_41_15_lpi_1;
  reg [11:0] buffer_bank3_data_41_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_41_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_21_14_12_lpi_1;
  reg buffer_bank3_data_21_15_lpi_1;
  reg [11:0] buffer_bank3_data_21_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_21_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_42_14_12_lpi_1;
  reg buffer_bank3_data_42_15_lpi_1;
  reg [11:0] buffer_bank3_data_42_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_42_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_20_14_12_lpi_1;
  reg buffer_bank3_data_20_15_lpi_1;
  reg [11:0] buffer_bank3_data_20_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_20_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_43_14_12_lpi_1;
  reg buffer_bank3_data_43_15_lpi_1;
  reg [11:0] buffer_bank3_data_43_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_43_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_19_14_12_lpi_1;
  reg buffer_bank3_data_19_15_lpi_1;
  reg [11:0] buffer_bank3_data_19_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_19_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_44_14_12_lpi_1;
  reg buffer_bank3_data_44_15_lpi_1;
  reg [11:0] buffer_bank3_data_44_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_44_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_18_14_12_lpi_1;
  reg buffer_bank3_data_18_15_lpi_1;
  reg [11:0] buffer_bank3_data_18_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_18_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_45_14_12_lpi_1;
  reg buffer_bank3_data_45_15_lpi_1;
  reg [11:0] buffer_bank3_data_45_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_45_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_17_14_12_lpi_1;
  reg buffer_bank3_data_17_15_lpi_1;
  reg [11:0] buffer_bank3_data_17_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_17_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_46_14_12_lpi_1;
  reg buffer_bank3_data_46_15_lpi_1;
  reg [11:0] buffer_bank3_data_46_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_46_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_16_14_12_lpi_1;
  reg buffer_bank3_data_16_15_lpi_1;
  reg [11:0] buffer_bank3_data_16_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_16_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_47_14_12_lpi_1;
  reg buffer_bank3_data_47_15_lpi_1;
  reg [11:0] buffer_bank3_data_47_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_47_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_15_14_12_lpi_1;
  reg buffer_bank3_data_15_15_lpi_1;
  reg [11:0] buffer_bank3_data_15_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_15_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_48_14_12_lpi_1;
  reg buffer_bank3_data_48_15_lpi_1;
  reg [11:0] buffer_bank3_data_48_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_48_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_14_14_12_lpi_1;
  reg buffer_bank3_data_14_15_lpi_1;
  reg [11:0] buffer_bank3_data_14_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_14_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_49_14_12_lpi_1;
  reg buffer_bank3_data_49_15_lpi_1;
  reg [11:0] buffer_bank3_data_49_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_49_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_13_14_12_lpi_1;
  reg buffer_bank3_data_13_15_lpi_1;
  reg [11:0] buffer_bank3_data_13_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_13_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_50_14_12_lpi_1;
  reg buffer_bank3_data_50_15_lpi_1;
  reg [11:0] buffer_bank3_data_50_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_50_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_12_14_12_lpi_1;
  reg buffer_bank3_data_12_15_lpi_1;
  reg [11:0] buffer_bank3_data_12_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_12_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_51_14_12_lpi_1;
  reg buffer_bank3_data_51_15_lpi_1;
  reg [11:0] buffer_bank3_data_51_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_51_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_11_14_12_lpi_1;
  reg buffer_bank3_data_11_15_lpi_1;
  reg [11:0] buffer_bank3_data_11_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_11_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_52_14_12_lpi_1;
  reg buffer_bank3_data_52_15_lpi_1;
  reg [11:0] buffer_bank3_data_52_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_52_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_10_14_12_lpi_1;
  reg buffer_bank3_data_10_15_lpi_1;
  reg [11:0] buffer_bank3_data_10_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_10_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_53_14_12_lpi_1;
  reg buffer_bank3_data_53_15_lpi_1;
  reg [11:0] buffer_bank3_data_53_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_53_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_9_14_12_lpi_1;
  reg buffer_bank3_data_9_15_lpi_1;
  reg [11:0] buffer_bank3_data_9_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_9_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_54_14_12_lpi_1;
  reg buffer_bank3_data_54_15_lpi_1;
  reg [11:0] buffer_bank3_data_54_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_54_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_8_14_12_lpi_1;
  reg buffer_bank3_data_8_15_lpi_1;
  reg [11:0] buffer_bank3_data_8_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_8_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_55_14_12_lpi_1;
  reg buffer_bank3_data_55_15_lpi_1;
  reg [11:0] buffer_bank3_data_55_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_55_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_7_14_12_lpi_1;
  reg buffer_bank3_data_7_15_lpi_1;
  reg [11:0] buffer_bank3_data_7_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_7_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_56_14_12_lpi_1;
  reg buffer_bank3_data_56_15_lpi_1;
  reg [11:0] buffer_bank3_data_56_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_56_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_6_14_12_lpi_1;
  reg buffer_bank3_data_6_15_lpi_1;
  reg [11:0] buffer_bank3_data_6_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_6_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_57_14_12_lpi_1;
  reg buffer_bank3_data_57_15_lpi_1;
  reg [11:0] buffer_bank3_data_57_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_57_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_5_14_12_lpi_1;
  reg buffer_bank3_data_5_15_lpi_1;
  reg [11:0] buffer_bank3_data_5_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_5_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_58_14_12_lpi_1;
  reg buffer_bank3_data_58_15_lpi_1;
  reg [11:0] buffer_bank3_data_58_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_58_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_4_14_12_lpi_1;
  reg buffer_bank3_data_4_15_lpi_1;
  reg [11:0] buffer_bank3_data_4_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_4_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_59_14_12_lpi_1;
  reg buffer_bank3_data_59_15_lpi_1;
  reg [11:0] buffer_bank3_data_59_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_59_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_3_14_12_lpi_1;
  reg buffer_bank3_data_3_15_lpi_1;
  reg [11:0] buffer_bank3_data_3_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_3_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_60_14_12_lpi_1;
  reg buffer_bank3_data_60_15_lpi_1;
  reg [11:0] buffer_bank3_data_60_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_60_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_2_14_12_lpi_1;
  reg buffer_bank3_data_2_15_lpi_1;
  reg [11:0] buffer_bank3_data_2_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_2_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_61_14_12_lpi_1;
  reg buffer_bank3_data_61_15_lpi_1;
  reg [11:0] buffer_bank3_data_61_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_61_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_1_14_12_lpi_1;
  reg buffer_bank3_data_1_15_lpi_1;
  reg [11:0] buffer_bank3_data_1_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_1_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_62_14_12_lpi_1;
  reg buffer_bank3_data_62_15_lpi_1;
  reg [11:0] buffer_bank3_data_62_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_62_31_16_lpi_1;
  reg [2:0] buffer_bank3_data_0_14_12_lpi_1;
  reg buffer_bank3_data_0_15_lpi_1;
  reg [11:0] buffer_bank3_data_0_11_0_lpi_1;
  reg [15:0] buffer_bank3_data_0_31_16_lpi_1;
  reg [9:0] buffer_bank4_data_31_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_31_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_32_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_32_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_30_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_30_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_33_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_33_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_29_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_29_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_34_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_34_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_28_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_28_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_35_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_35_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_27_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_27_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_36_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_36_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_26_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_26_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_37_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_37_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_25_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_25_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_38_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_38_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_24_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_24_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_39_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_39_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_23_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_23_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_40_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_40_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_22_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_22_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_41_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_41_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_21_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_21_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_42_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_42_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_20_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_20_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_43_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_43_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_19_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_19_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_44_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_44_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_18_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_18_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_45_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_45_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_17_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_17_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_46_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_46_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_16_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_16_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_47_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_47_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_15_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_15_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_48_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_48_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_14_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_14_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_49_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_49_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_13_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_13_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_50_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_50_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_12_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_12_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_51_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_51_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_11_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_11_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_52_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_52_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_10_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_10_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_53_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_53_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_9_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_9_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_54_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_54_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_8_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_8_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_55_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_55_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_7_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_7_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_56_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_56_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_6_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_6_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_57_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_57_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_5_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_5_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_58_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_58_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_4_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_4_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_59_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_59_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_3_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_3_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_60_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_60_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_2_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_2_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_61_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_61_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_1_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_1_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_62_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_62_31_10_lpi_1;
  reg [9:0] buffer_bank4_data_0_9_0_lpi_1;
  reg [21:0] buffer_bank4_data_0_31_10_lpi_1;
  reg [25:0] buffer_bank5_data_31_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_31_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_31_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_32_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_32_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_32_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_30_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_30_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_30_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_33_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_33_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_33_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_29_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_29_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_29_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_34_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_34_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_34_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_28_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_28_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_28_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_35_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_35_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_35_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_27_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_27_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_27_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_36_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_36_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_36_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_26_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_26_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_26_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_37_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_37_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_37_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_25_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_25_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_25_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_38_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_38_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_38_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_24_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_24_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_24_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_39_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_39_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_39_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_23_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_23_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_23_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_40_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_40_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_40_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_22_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_22_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_22_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_41_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_41_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_41_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_21_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_21_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_21_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_42_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_42_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_42_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_20_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_20_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_20_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_43_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_43_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_43_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_19_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_19_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_19_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_44_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_44_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_44_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_18_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_18_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_18_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_45_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_45_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_45_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_17_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_17_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_17_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_46_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_46_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_46_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_16_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_16_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_16_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_47_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_47_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_47_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_15_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_15_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_15_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_48_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_48_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_48_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_14_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_14_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_14_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_49_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_49_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_49_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_13_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_13_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_13_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_50_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_50_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_50_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_12_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_12_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_12_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_51_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_51_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_51_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_11_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_11_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_11_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_52_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_52_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_52_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_10_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_10_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_10_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_53_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_53_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_53_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_9_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_9_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_9_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_54_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_54_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_54_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_8_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_8_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_8_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_55_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_55_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_55_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_7_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_7_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_7_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_56_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_56_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_56_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_6_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_6_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_6_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_57_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_57_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_57_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_5_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_5_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_5_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_58_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_58_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_58_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_4_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_4_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_4_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_59_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_59_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_59_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_3_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_3_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_3_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_60_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_60_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_60_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_2_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_2_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_2_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_61_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_61_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_61_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_1_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_1_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_1_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_62_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_62_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_62_31_30_lpi_1;
  reg [25:0] buffer_bank5_data_0_29_4_lpi_1;
  reg [3:0] buffer_bank5_data_0_3_0_lpi_1;
  reg [1:0] buffer_bank5_data_0_31_30_lpi_1;
  reg [22:0] buffer_bank6_data_31_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_31_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_32_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_32_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_30_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_30_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_33_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_33_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_29_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_29_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_34_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_34_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_28_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_28_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_35_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_35_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_27_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_27_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_36_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_36_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_26_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_26_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_37_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_37_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_25_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_25_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_38_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_38_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_24_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_24_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_39_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_39_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_23_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_23_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_40_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_40_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_22_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_22_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_41_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_41_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_21_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_21_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_42_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_42_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_20_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_20_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_43_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_43_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_19_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_19_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_44_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_44_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_18_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_18_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_45_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_45_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_17_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_17_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_46_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_46_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_16_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_16_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_47_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_47_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_15_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_15_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_48_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_48_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_14_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_14_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_49_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_49_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_13_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_13_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_50_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_50_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_12_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_12_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_51_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_51_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_11_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_11_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_52_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_52_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_10_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_10_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_53_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_53_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_9_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_9_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_54_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_54_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_8_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_8_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_55_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_55_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_7_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_7_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_56_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_56_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_6_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_6_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_57_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_57_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_5_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_5_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_58_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_58_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_4_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_4_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_59_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_59_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_3_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_3_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_60_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_60_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_2_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_2_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_61_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_61_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_1_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_1_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_62_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_62_31_23_lpi_1;
  reg [22:0] buffer_bank6_data_0_22_0_lpi_1;
  reg [8:0] buffer_bank6_data_0_31_23_lpi_1;
  reg [15:0] buffer_bank7_data_31_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_31_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_32_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_32_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_30_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_30_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_33_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_33_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_29_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_29_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_34_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_34_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_28_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_28_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_35_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_35_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_27_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_27_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_36_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_36_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_26_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_26_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_37_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_37_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_25_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_25_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_38_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_38_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_24_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_24_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_39_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_39_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_23_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_23_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_40_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_40_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_22_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_22_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_41_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_41_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_21_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_21_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_42_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_42_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_20_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_20_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_43_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_43_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_19_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_19_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_44_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_44_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_18_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_18_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_45_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_45_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_17_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_17_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_46_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_46_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_16_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_16_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_47_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_47_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_15_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_15_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_48_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_48_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_14_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_14_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_49_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_49_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_13_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_13_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_50_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_50_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_12_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_12_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_51_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_51_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_11_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_11_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_52_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_52_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_10_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_10_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_53_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_53_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_9_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_9_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_54_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_54_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_8_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_8_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_55_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_55_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_7_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_7_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_56_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_56_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_6_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_6_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_57_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_57_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_5_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_5_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_58_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_58_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_4_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_4_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_59_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_59_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_3_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_3_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_60_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_60_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_2_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_2_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_61_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_61_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_1_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_1_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_62_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_62_31_16_lpi_1;
  reg [15:0] buffer_bank7_data_0_15_0_lpi_1;
  reg [15:0] buffer_bank7_data_0_31_16_lpi_1;
  reg [8:0] buffer_bank8_data_31_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_31_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_32_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_32_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_30_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_30_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_33_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_33_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_29_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_29_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_34_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_34_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_28_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_28_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_35_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_35_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_27_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_27_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_36_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_36_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_26_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_26_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_37_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_37_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_25_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_25_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_38_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_38_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_24_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_24_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_39_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_39_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_23_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_23_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_40_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_40_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_22_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_22_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_41_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_41_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_21_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_21_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_42_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_42_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_20_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_20_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_43_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_43_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_19_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_19_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_44_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_44_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_18_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_18_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_45_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_45_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_17_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_17_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_46_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_46_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_16_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_16_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_47_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_47_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_15_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_15_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_48_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_48_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_14_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_14_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_49_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_49_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_13_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_13_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_50_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_50_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_12_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_12_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_51_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_51_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_11_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_11_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_52_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_52_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_10_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_10_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_53_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_53_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_9_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_9_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_54_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_54_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_8_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_8_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_55_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_55_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_7_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_7_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_56_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_56_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_6_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_6_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_57_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_57_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_5_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_5_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_58_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_58_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_4_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_4_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_59_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_59_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_3_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_3_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_60_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_60_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_2_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_2_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_61_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_61_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_1_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_1_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_62_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_62_31_9_lpi_1;
  reg [8:0] buffer_bank8_data_0_8_0_lpi_1;
  reg [22:0] buffer_bank8_data_0_31_9_lpi_1;
  reg [7:0] buffer_bank9_data_31_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_31_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_32_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_32_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_30_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_30_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_33_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_33_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_29_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_29_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_34_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_34_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_28_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_28_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_35_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_35_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_27_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_27_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_36_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_36_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_26_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_26_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_37_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_37_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_25_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_25_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_38_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_38_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_24_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_24_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_39_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_39_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_23_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_23_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_40_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_40_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_22_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_22_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_41_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_41_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_21_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_21_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_42_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_42_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_20_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_20_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_43_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_43_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_19_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_19_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_44_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_44_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_18_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_18_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_45_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_45_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_17_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_17_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_46_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_46_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_16_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_16_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_47_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_47_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_15_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_15_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_48_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_48_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_14_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_14_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_49_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_49_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_13_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_13_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_50_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_50_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_12_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_12_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_51_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_51_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_11_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_11_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_52_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_52_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_10_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_10_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_53_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_53_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_9_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_9_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_54_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_54_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_8_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_8_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_55_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_55_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_7_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_7_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_56_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_56_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_6_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_6_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_57_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_57_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_5_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_5_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_58_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_58_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_4_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_4_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_59_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_59_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_3_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_3_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_60_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_60_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_2_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_2_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_61_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_61_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_1_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_1_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_62_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_62_31_8_lpi_1;
  reg [7:0] buffer_bank9_data_0_7_0_lpi_1;
  reg [23:0] buffer_bank9_data_0_31_8_lpi_1;
  reg [26:0] buffer_bank10_data_31_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_31_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_31_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_32_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_32_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_32_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_30_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_30_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_30_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_33_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_33_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_33_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_29_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_29_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_29_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_34_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_34_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_34_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_28_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_28_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_28_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_35_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_35_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_35_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_27_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_27_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_27_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_36_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_36_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_36_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_26_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_26_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_26_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_37_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_37_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_37_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_25_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_25_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_25_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_38_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_38_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_38_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_24_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_24_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_24_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_39_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_39_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_39_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_23_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_23_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_23_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_40_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_40_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_40_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_22_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_22_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_22_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_41_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_41_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_41_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_21_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_21_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_21_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_42_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_42_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_42_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_20_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_20_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_20_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_43_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_43_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_43_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_19_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_19_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_19_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_44_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_44_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_44_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_18_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_18_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_18_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_45_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_45_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_45_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_17_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_17_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_17_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_46_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_46_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_46_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_16_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_16_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_16_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_47_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_47_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_47_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_15_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_15_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_15_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_48_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_48_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_48_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_14_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_14_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_14_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_49_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_49_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_49_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_13_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_13_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_13_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_50_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_50_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_50_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_12_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_12_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_12_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_51_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_51_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_51_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_11_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_11_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_11_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_52_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_52_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_52_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_10_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_10_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_10_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_53_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_53_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_53_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_9_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_9_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_9_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_54_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_54_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_54_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_8_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_8_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_8_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_55_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_55_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_55_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_7_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_7_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_7_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_56_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_56_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_56_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_6_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_6_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_6_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_57_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_57_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_57_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_5_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_5_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_5_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_58_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_58_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_58_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_4_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_4_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_4_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_59_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_59_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_59_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_3_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_3_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_3_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_60_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_60_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_60_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_2_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_2_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_2_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_61_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_61_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_61_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_1_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_1_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_1_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_62_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_62_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_62_31_30_lpi_1;
  reg [26:0] buffer_bank10_data_0_29_3_lpi_1;
  reg [2:0] buffer_bank10_data_0_2_0_lpi_1;
  reg [1:0] buffer_bank10_data_0_31_30_lpi_1;
  reg [24:0] buffer_bank11_data_31_lpi_1;
  reg [24:0] buffer_bank11_data_32_lpi_1;
  reg [24:0] buffer_bank11_data_30_lpi_1;
  reg [24:0] buffer_bank11_data_33_lpi_1;
  reg [24:0] buffer_bank11_data_29_lpi_1;
  reg [24:0] buffer_bank11_data_34_lpi_1;
  reg [24:0] buffer_bank11_data_28_lpi_1;
  reg [24:0] buffer_bank11_data_35_lpi_1;
  reg [24:0] buffer_bank11_data_27_lpi_1;
  reg [24:0] buffer_bank11_data_36_lpi_1;
  reg [24:0] buffer_bank11_data_26_lpi_1;
  reg [24:0] buffer_bank11_data_37_lpi_1;
  reg [24:0] buffer_bank11_data_25_lpi_1;
  reg [24:0] buffer_bank11_data_38_lpi_1;
  reg [24:0] buffer_bank11_data_24_lpi_1;
  reg [24:0] buffer_bank11_data_39_lpi_1;
  reg [24:0] buffer_bank11_data_23_lpi_1;
  reg [24:0] buffer_bank11_data_40_lpi_1;
  reg [24:0] buffer_bank11_data_22_lpi_1;
  reg [24:0] buffer_bank11_data_41_lpi_1;
  reg [24:0] buffer_bank11_data_21_lpi_1;
  reg [24:0] buffer_bank11_data_42_lpi_1;
  reg [24:0] buffer_bank11_data_20_lpi_1;
  reg [24:0] buffer_bank11_data_43_lpi_1;
  reg [24:0] buffer_bank11_data_19_lpi_1;
  reg [24:0] buffer_bank11_data_44_lpi_1;
  reg [24:0] buffer_bank11_data_18_lpi_1;
  reg [24:0] buffer_bank11_data_45_lpi_1;
  reg [24:0] buffer_bank11_data_17_lpi_1;
  reg [24:0] buffer_bank11_data_46_lpi_1;
  reg [24:0] buffer_bank11_data_16_lpi_1;
  reg [24:0] buffer_bank11_data_47_lpi_1;
  reg [24:0] buffer_bank11_data_15_lpi_1;
  reg [24:0] buffer_bank11_data_48_lpi_1;
  reg [24:0] buffer_bank11_data_14_lpi_1;
  reg [24:0] buffer_bank11_data_49_lpi_1;
  reg [24:0] buffer_bank11_data_13_lpi_1;
  reg [24:0] buffer_bank11_data_50_lpi_1;
  reg [24:0] buffer_bank11_data_12_lpi_1;
  reg [24:0] buffer_bank11_data_51_lpi_1;
  reg [24:0] buffer_bank11_data_11_lpi_1;
  reg [24:0] buffer_bank11_data_52_lpi_1;
  reg [24:0] buffer_bank11_data_10_lpi_1;
  reg [24:0] buffer_bank11_data_53_lpi_1;
  reg [24:0] buffer_bank11_data_9_lpi_1;
  reg [24:0] buffer_bank11_data_54_lpi_1;
  reg [24:0] buffer_bank11_data_8_lpi_1;
  reg [24:0] buffer_bank11_data_55_lpi_1;
  reg [24:0] buffer_bank11_data_7_lpi_1;
  reg [24:0] buffer_bank11_data_56_lpi_1;
  reg [24:0] buffer_bank11_data_6_lpi_1;
  reg [24:0] buffer_bank11_data_57_lpi_1;
  reg [24:0] buffer_bank11_data_5_lpi_1;
  reg [24:0] buffer_bank11_data_58_lpi_1;
  reg [24:0] buffer_bank11_data_4_lpi_1;
  reg [24:0] buffer_bank11_data_59_lpi_1;
  reg [24:0] buffer_bank11_data_3_lpi_1;
  reg [24:0] buffer_bank11_data_60_lpi_1;
  reg [24:0] buffer_bank11_data_2_lpi_1;
  reg [24:0] buffer_bank11_data_61_lpi_1;
  reg [24:0] buffer_bank11_data_1_lpi_1;
  reg [24:0] buffer_bank11_data_62_lpi_1;
  reg [24:0] buffer_bank11_data_0_lpi_1;
  reg [376:0] quads_in_crt_lpi_1;
  reg exit_for_sva;
  reg operator_2_false_2_operator_2_false_2_and_mdf_sva_1;
  reg operator_2_false_1_operator_2_false_1_and_mdf_sva_1;
  reg operator_2_false_operator_2_false_nor_mdf_sva_1;
  reg [5:0] for_1_for_quad_idx_lpi_1_5_0;
  reg [32:0] paramsIn_crt_lpi_1_dfm_56_24;
  reg [12:0] paramsIn_crt_lpi_1_dfm_12_0;
  wire [5:0] for_1_for_quad_idx_lpi_1_dfm_5_0_1;
  wire [32:0] paramsIn_crt_lpi_1_dfm_56_24_mx0;
  wire qelse_qelse_and_cse;
  wire for_and_123_cse;
  wire buffer_bank11_data_and_cse;
  wire buffer_bank11_data_and_1_cse;
  wire buffer_bank11_data_and_2_cse;
  wire buffer_bank11_data_and_3_cse;
  wire buffer_bank11_data_and_4_cse;
  wire buffer_bank11_data_and_5_cse;
  wire buffer_bank11_data_and_6_cse;
  wire buffer_bank11_data_and_7_cse;
  wire buffer_bank11_data_and_8_cse;
  wire buffer_bank11_data_and_9_cse;
  wire buffer_bank11_data_and_10_cse;
  wire buffer_bank11_data_and_11_cse;
  wire buffer_bank11_data_and_12_cse;
  wire buffer_bank11_data_and_13_cse;
  wire buffer_bank11_data_and_14_cse;
  wire buffer_bank11_data_and_15_cse;
  wire buffer_bank11_data_and_16_cse;
  wire buffer_bank11_data_and_17_cse;
  wire buffer_bank11_data_and_18_cse;
  wire buffer_bank11_data_and_19_cse;
  wire buffer_bank11_data_and_20_cse;
  wire buffer_bank11_data_and_21_cse;
  wire buffer_bank11_data_and_22_cse;
  wire buffer_bank11_data_and_23_cse;
  wire buffer_bank11_data_and_24_cse;
  wire buffer_bank11_data_and_25_cse;
  wire buffer_bank11_data_and_26_cse;
  wire buffer_bank11_data_and_27_cse;
  wire buffer_bank11_data_and_28_cse;
  wire buffer_bank11_data_and_29_cse;
  wire buffer_bank11_data_and_30_cse;
  wire buffer_bank11_data_and_31_cse;
  wire buffer_bank11_data_and_32_cse;
  wire buffer_bank11_data_and_33_cse;
  wire buffer_bank11_data_and_34_cse;
  wire buffer_bank11_data_and_35_cse;
  wire buffer_bank11_data_and_36_cse;
  wire buffer_bank11_data_and_37_cse;
  wire buffer_bank11_data_and_38_cse;
  wire buffer_bank11_data_and_39_cse;
  wire buffer_bank11_data_and_40_cse;
  wire buffer_bank11_data_and_41_cse;
  wire buffer_bank11_data_and_42_cse;
  wire buffer_bank11_data_and_43_cse;
  wire buffer_bank11_data_and_44_cse;
  wire buffer_bank11_data_and_45_cse;
  wire buffer_bank11_data_and_46_cse;
  wire buffer_bank11_data_and_47_cse;
  wire buffer_bank11_data_and_48_cse;
  wire buffer_bank11_data_and_49_cse;
  wire buffer_bank11_data_and_50_cse;
  wire buffer_bank11_data_and_51_cse;
  wire buffer_bank11_data_and_52_cse;
  wire buffer_bank11_data_and_53_cse;
  wire buffer_bank11_data_and_54_cse;
  wire buffer_bank11_data_and_55_cse;
  wire buffer_bank11_data_and_56_cse;
  wire buffer_bank11_data_and_57_cse;
  wire buffer_bank11_data_and_58_cse;
  wire buffer_bank11_data_and_59_cse;
  wire buffer_bank11_data_and_60_cse;
  wire buffer_bank11_data_and_61_cse;
  wire buffer_bank11_data_and_62_cse;
  wire for_1_if_equal_tmp;
  wire mux_tmp_89;
  wire mux_tmp_91;
  wire mux_tmp_93;
  wire nor_tmp_14;
  wire or_tmp_183;
  wire and_tmp_2;
  wire nor_tmp_15;
  wire and_tmp_3;
  wire for_1_and_1901_cse;
  wire or_1_cse;
  wire or_297_cse;
  wire or_302_cse;
  wire operator_43_false_acc_itm_43;

  wire[21:0] pixels_in_img_mul_nl;
  wire signed [23:0] nl_pixels_in_img_mul_nl;
  wire[0:0] nor_30_nl;
  wire[0:0] for_1_not_3868_nl;
  wire[0:0] mux_93_nl;
  wire[0:0] nor_100_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_97_nl;
  wire[0:0] or_303_nl;
  wire[0:0] nand_12_nl;
  wire[42:0] for_for_and_nl;
  wire[0:0] for_1_for_1_for_not_1_nl;
  wire[0:0] for_1_and_1900_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] mux_102_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] or_300_nl;
  wire[0:0] or_299_nl;
  wire[0:0] mux_101_nl;
  wire[0:0] mux_100_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] nand_10_nl;
  wire[0:0] or_298_nl;
  wire[0:0] mux_98_nl;
  wire[0:0] or_292_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] or_15_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_13_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] or_11_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] or_9_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nand_8_nl;
  wire[0:0] or_164_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] for_for_or_nl;
  wire[0:0] nor_nl;
  wire[0:0] and_1_nl;
  wire[0:0] and_2_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] for_1_mux_1960_nl;
  wire[0:0] for_1_for_mux_5_nl;
  wire[0:0] for_1_and_1893_nl;
  wire[0:0] for_1_and_1894_nl;
  wire[0:0] and_32_nl;
  wire[10:0] for_1_mux_3_nl;
  wire[24:0] for_1_mux_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] for_1_not_3876_nl;
  wire[0:0] for_1_for_1_for_nor_nl;
  wire[43:0] operator_43_false_acc_nl;
  wire[44:0] nl_operator_43_false_acc_nl;
  wire[0:0] or_279_nl;
  wire[0:0] for_1_for_1_nor_1894_nl;
  wire[0:0] for_mux_nl;
  wire[0:0] or_8_nl;
  wire[0:0] or_7_nl;
  wire[0:0] or_19_nl;
  wire[0:0] or_22_nl;
  wire[0:0] or_24_nl;
  wire[0:0] or_26_nl;
  wire[0:0] or_28_nl;
  wire[0:0] or_30_nl;
  wire[0:0] or_32_nl;
  wire[0:0] or_34_nl;
  wire[0:0] or_36_nl;
  wire[0:0] or_38_nl;
  wire[0:0] or_40_nl;
  wire[0:0] or_42_nl;
  wire[0:0] or_44_nl;
  wire[0:0] or_46_nl;
  wire[0:0] or_48_nl;
  wire[0:0] or_50_nl;
  wire[0:0] or_52_nl;
  wire[0:0] or_54_nl;
  wire[0:0] or_56_nl;
  wire[0:0] or_58_nl;
  wire[0:0] or_60_nl;
  wire[0:0] or_62_nl;
  wire[0:0] or_64_nl;
  wire[0:0] or_66_nl;
  wire[0:0] or_68_nl;
  wire[0:0] or_70_nl;
  wire[0:0] or_72_nl;
  wire[0:0] or_74_nl;
  wire[0:0] or_76_nl;
  wire[0:0] or_78_nl;
  wire[0:0] or_80_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] or_84_nl;
  wire[0:0] or_86_nl;
  wire[0:0] or_88_nl;
  wire[0:0] or_90_nl;
  wire[0:0] or_92_nl;
  wire[0:0] or_94_nl;
  wire[0:0] or_96_nl;
  wire[0:0] or_98_nl;
  wire[0:0] or_100_nl;
  wire[0:0] or_102_nl;
  wire[0:0] or_104_nl;
  wire[0:0] or_106_nl;
  wire[0:0] or_108_nl;
  wire[0:0] or_110_nl;
  wire[0:0] or_112_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] or_116_nl;
  wire[0:0] or_118_nl;
  wire[0:0] or_120_nl;
  wire[0:0] or_122_nl;
  wire[0:0] or_124_nl;
  wire[0:0] or_126_nl;
  wire[0:0] or_128_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] or_132_nl;
  wire[0:0] or_134_nl;
  wire[0:0] or_136_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] or_140_nl;
  wire[0:0] nand_5_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] or_287_nl;
  wire[0:0] or_286_nl;
  wire[0:0] or_289_nl;
  wire[0:0] mux_95_nl;
  wire[0:0] or_288_nl;
  wire[0:0] and_38_nl;
  wire[43:0] acc_nl;
  wire[44:0] nl_acc_nl;
  wire[42:0] pixels_in_img_mux_2_nl;
  wire[10:0] pixels_in_img_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [376:0] nl_QuadBuffer_64_run_quads_out_rsci_inst_quads_out_rsci_idat;
  assign nl_QuadBuffer_64_run_quads_out_rsci_inst_quads_out_rsci_idat = {quads_out_rsci_idat_376_352
      , quads_out_rsci_idat_351_350 , quads_out_rsci_idat_349_323 , quads_out_rsci_idat_322_320
      , quads_out_rsci_idat_319_296 , quads_out_rsci_idat_295_288 , quads_out_rsci_idat_287_265
      , quads_out_rsci_idat_264_256 , quads_out_rsci_idat_255_240 , quads_out_rsci_idat_239_224
      , quads_out_rsci_idat_223_215 , quads_out_rsci_idat_214_192 , quads_out_rsci_idat_191_190
      , quads_out_rsci_idat_189_164 , quads_out_rsci_idat_163_160 , quads_out_rsci_idat_159_138
      , quads_out_rsci_idat_137_128 , quads_out_rsci_idat_127_112 , quads_out_rsci_idat_111
      , quads_out_rsci_idat_110_108 , quads_out_rsci_idat_107_96 , quads_out_rsci_idat_95_84
      , quads_out_rsci_idat_83_72 , quads_out_rsci_idat_71_64 , quads_out_rsci_idat_63_60
      , quads_out_rsci_idat_59_48 , quads_out_rsci_idat_47_36 , quads_out_rsci_idat_35_32
      , quads_out_rsci_idat_31_24 , quads_out_rsci_idat_23_12 , quads_out_rsci_idat_11_0};
  QuadBuffer_64_run_quads_in_rsci QuadBuffer_64_run_quads_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsc_dat(quads_in_rsc_dat),
      .quads_in_rsc_vld(quads_in_rsc_vld),
      .quads_in_rsc_rdy(quads_in_rsc_rdy),
      .run_wen(run_wen),
      .quads_in_rsci_oswt(reg_quads_in_rsci_oswt_cse),
      .quads_in_rsci_wen_comp(quads_in_rsci_wen_comp),
      .quads_in_rsci_idat_mxwt(quads_in_rsci_idat_mxwt)
    );
  QuadBuffer_64_run_paramsIn_rsci QuadBuffer_64_run_paramsIn_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_oswt_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  QuadBuffer_64_run_quads_out_rsci QuadBuffer_64_run_quads_out_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_out_rsc_dat(quads_out_rsc_dat),
      .quads_out_rsc_vld(quads_out_rsc_vld),
      .quads_out_rsc_rdy(quads_out_rsc_rdy),
      .run_wen(run_wen),
      .quads_out_rsci_oswt(reg_quads_out_rsci_oswt_cse),
      .quads_out_rsci_wen_comp(quads_out_rsci_wen_comp),
      .quads_out_rsci_idat(nl_QuadBuffer_64_run_quads_out_rsci_inst_quads_out_rsci_idat[376:0])
    );
  QuadBuffer_64_run_staller QuadBuffer_64_run_staller_inst (
      .run_wen(run_wen),
      .quads_in_rsci_wen_comp(quads_in_rsci_wen_comp),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .quads_out_rsci_wen_comp(quads_out_rsci_wen_comp)
    );
  assign qelse_qelse_and_cse = run_wen & and_dcpl_7;
  assign quads_out_and_cse = run_wen & (~ or_dcpl_13);
  assign nor_30_nl = ~((for_1_mux1h_2098_tmp!=2'b00));
  assign mux_89_cse = MUX_s_1_2_2(exitL_exit_for_1_sva, (nor_30_nl), main_stage_0_2);
  assign or_1_cse = (for_1_mux1h_2098_tmp!=2'b00);
  assign mux_4_nl = MUX_s_1_2_2((~ exitL_exit_for_1_sva), (for_1_mux1h_2098_tmp[1]),
      main_stage_0_2);
  assign for_and_123_cse = run_wen & (mux_4_nl) & (~ or_dcpl_2);
  assign or_297_cse = (operator_11_false_2_acc_tmp[11:6]!=6'b000000);
  assign buffer_bank11_data_and_cse = run_wen & mux_tmp_9 & (~(or_dcpl_18 | or_dcpl_16));
  assign buffer_bank11_data_and_1_cse = run_wen & mux_tmp_10 & (~(or_dcpl_21 | or_dcpl_16));
  assign buffer_bank11_data_and_2_cse = run_wen & mux_tmp_11 & (~(or_dcpl_24 | or_dcpl_16));
  assign buffer_bank11_data_and_3_cse = run_wen & mux_tmp_12 & (~(or_dcpl_27 | or_dcpl_16));
  assign buffer_bank11_data_and_4_cse = run_wen & mux_tmp_13 & (~(or_dcpl_18 | or_dcpl_30));
  assign buffer_bank11_data_and_5_cse = run_wen & mux_tmp_14 & (~(or_dcpl_21 | or_dcpl_30));
  assign buffer_bank11_data_and_6_cse = run_wen & mux_tmp_15 & (~(or_dcpl_24 | or_dcpl_30));
  assign buffer_bank11_data_and_7_cse = run_wen & mux_tmp_16 & (~(or_dcpl_27 | or_dcpl_30));
  assign buffer_bank11_data_and_8_cse = run_wen & mux_tmp_17 & (~(or_dcpl_18 | or_dcpl_36));
  assign buffer_bank11_data_and_9_cse = run_wen & mux_tmp_18 & (~(or_dcpl_21 | or_dcpl_36));
  assign buffer_bank11_data_and_10_cse = run_wen & mux_tmp_19 & (~(or_dcpl_24 | or_dcpl_36));
  assign buffer_bank11_data_and_11_cse = run_wen & mux_tmp_20 & (~(or_dcpl_27 | or_dcpl_36));
  assign buffer_bank11_data_and_12_cse = run_wen & mux_tmp_21 & (~(or_dcpl_18 | or_dcpl_42));
  assign buffer_bank11_data_and_13_cse = run_wen & mux_tmp_22 & (~(or_dcpl_21 | or_dcpl_42));
  assign buffer_bank11_data_and_14_cse = run_wen & mux_tmp_23 & (~(or_dcpl_24 | or_dcpl_42));
  assign buffer_bank11_data_and_15_cse = run_wen & mux_tmp_24 & (~(or_dcpl_27 | or_dcpl_42));
  assign buffer_bank11_data_and_16_cse = run_wen & mux_tmp_25 & (~(or_dcpl_18 | or_dcpl_48));
  assign buffer_bank11_data_and_17_cse = run_wen & mux_tmp_26 & (~(or_dcpl_21 | or_dcpl_48));
  assign buffer_bank11_data_and_18_cse = run_wen & mux_tmp_27 & (~(or_dcpl_24 | or_dcpl_48));
  assign buffer_bank11_data_and_19_cse = run_wen & mux_tmp_28 & (~(or_dcpl_27 | or_dcpl_48));
  assign buffer_bank11_data_and_20_cse = run_wen & mux_tmp_29 & (~(or_dcpl_18 | or_dcpl_53));
  assign buffer_bank11_data_and_21_cse = run_wen & mux_tmp_30 & (~(or_dcpl_21 | or_dcpl_53));
  assign buffer_bank11_data_and_22_cse = run_wen & mux_tmp_31 & (~(or_dcpl_24 | or_dcpl_53));
  assign buffer_bank11_data_and_23_cse = run_wen & mux_tmp_32 & (~(or_dcpl_27 | or_dcpl_53));
  assign buffer_bank11_data_and_24_cse = run_wen & mux_tmp_33 & (~(or_dcpl_18 | or_dcpl_58));
  assign buffer_bank11_data_and_25_cse = run_wen & mux_tmp_34 & (~(or_dcpl_21 | or_dcpl_58));
  assign buffer_bank11_data_and_26_cse = run_wen & mux_tmp_35 & (~(or_dcpl_24 | or_dcpl_58));
  assign buffer_bank11_data_and_27_cse = run_wen & mux_tmp_36 & (~(or_dcpl_27 | or_dcpl_58));
  assign buffer_bank11_data_and_28_cse = run_wen & mux_tmp_37 & (~(or_dcpl_18 | or_dcpl_63));
  assign buffer_bank11_data_and_29_cse = run_wen & mux_tmp_38 & (~(or_dcpl_21 | or_dcpl_63));
  assign buffer_bank11_data_and_30_cse = run_wen & mux_tmp_39 & (~(or_dcpl_24 | or_dcpl_63));
  assign buffer_bank11_data_and_31_cse = run_wen & mux_tmp_40 & (~(or_dcpl_27 | or_dcpl_63));
  assign buffer_bank11_data_and_32_cse = run_wen & mux_tmp_41 & (~(or_dcpl_18 | or_dcpl_69));
  assign buffer_bank11_data_and_33_cse = run_wen & mux_tmp_42 & (~(or_dcpl_21 | or_dcpl_69));
  assign buffer_bank11_data_and_34_cse = run_wen & mux_tmp_43 & (~(or_dcpl_24 | or_dcpl_69));
  assign buffer_bank11_data_and_35_cse = run_wen & mux_tmp_44 & (~(or_dcpl_27 | or_dcpl_69));
  assign buffer_bank11_data_and_36_cse = run_wen & mux_tmp_45 & (~(or_dcpl_18 | or_dcpl_74));
  assign buffer_bank11_data_and_37_cse = run_wen & mux_tmp_46 & (~(or_dcpl_21 | or_dcpl_74));
  assign buffer_bank11_data_and_38_cse = run_wen & mux_tmp_47 & (~(or_dcpl_24 | or_dcpl_74));
  assign buffer_bank11_data_and_39_cse = run_wen & mux_tmp_48 & (~(or_dcpl_27 | or_dcpl_74));
  assign buffer_bank11_data_and_40_cse = run_wen & mux_tmp_49 & (~(or_dcpl_18 | or_dcpl_79));
  assign buffer_bank11_data_and_41_cse = run_wen & mux_tmp_50 & (~(or_dcpl_21 | or_dcpl_79));
  assign buffer_bank11_data_and_42_cse = run_wen & mux_tmp_51 & (~(or_dcpl_24 | or_dcpl_79));
  assign buffer_bank11_data_and_43_cse = run_wen & mux_tmp_52 & (~(or_dcpl_27 | or_dcpl_79));
  assign buffer_bank11_data_and_44_cse = run_wen & mux_tmp_53 & (~(or_dcpl_18 | or_dcpl_84));
  assign buffer_bank11_data_and_45_cse = run_wen & mux_tmp_54 & (~(or_dcpl_21 | or_dcpl_84));
  assign buffer_bank11_data_and_46_cse = run_wen & mux_tmp_55 & (~(or_dcpl_24 | or_dcpl_84));
  assign buffer_bank11_data_and_47_cse = run_wen & mux_tmp_56 & (~(or_dcpl_27 | or_dcpl_84));
  assign buffer_bank11_data_and_48_cse = run_wen & mux_tmp_57 & (~(or_dcpl_18 | or_dcpl_90));
  assign buffer_bank11_data_and_49_cse = run_wen & mux_tmp_58 & (~(or_dcpl_21 | or_dcpl_90));
  assign buffer_bank11_data_and_50_cse = run_wen & mux_tmp_59 & (~(or_dcpl_24 | or_dcpl_90));
  assign buffer_bank11_data_and_51_cse = run_wen & mux_tmp_60 & (~(or_dcpl_27 | or_dcpl_90));
  assign buffer_bank11_data_and_52_cse = run_wen & mux_tmp_61 & (~(or_dcpl_18 | or_dcpl_95));
  assign buffer_bank11_data_and_53_cse = run_wen & mux_tmp_62 & (~(or_dcpl_21 | or_dcpl_95));
  assign buffer_bank11_data_and_54_cse = run_wen & mux_tmp_63 & (~(or_dcpl_24 | or_dcpl_95));
  assign buffer_bank11_data_and_55_cse = run_wen & mux_tmp_64 & (~(or_dcpl_27 | or_dcpl_95));
  assign buffer_bank11_data_and_56_cse = run_wen & mux_tmp_65 & (~(or_dcpl_18 | or_dcpl_100));
  assign buffer_bank11_data_and_57_cse = run_wen & mux_tmp_66 & (~(or_dcpl_21 | or_dcpl_100));
  assign buffer_bank11_data_and_58_cse = run_wen & mux_tmp_67 & (~(or_dcpl_24 | or_dcpl_100));
  assign buffer_bank11_data_and_59_cse = run_wen & mux_tmp_68 & (~(or_dcpl_27 | or_dcpl_100));
  assign buffer_bank11_data_and_60_cse = run_wen & mux_tmp_69 & (~(or_dcpl_18 | or_dcpl_105));
  assign buffer_bank11_data_and_61_cse = run_wen & mux_tmp_70 & (~(or_dcpl_21 | or_dcpl_105));
  assign buffer_bank11_data_and_62_cse = run_wen & mux_tmp_71 & (~(or_dcpl_24 | or_dcpl_105));
  assign for_1_and_1901_cse = run_wen & main_stage_0_2;
  assign nor_nl = ~(operator_2_false_2_operator_2_false_2_and_mdf_sva_1 | operator_2_false_1_operator_2_false_1_and_mdf_sva_1
      | operator_2_false_operator_2_false_nor_mdf_sva_1);
  assign and_1_nl = operator_2_false_2_operator_2_false_2_and_mdf_sva_1 & (~ operator_2_false_1_operator_2_false_1_and_mdf_sva_1)
      & (~ operator_2_false_operator_2_false_nor_mdf_sva_1);
  assign and_2_nl = operator_2_false_1_operator_2_false_1_and_mdf_sva_1 & (~ operator_2_false_operator_2_false_nor_mdf_sva_1);
  assign nl_tot_samples_in_img_mul_psp_sva_1 = (tot_samples_in_img_mul_psp_lpi_1[21:0])
      * ({(nor_nl) , 1'b0 , (and_1_nl) , 1'b0 , (and_2_nl) , operator_2_false_operator_2_false_nor_mdf_sva_1});
  assign tot_samples_in_img_mul_psp_sva_1 = nl_tot_samples_in_img_mul_psp_sva_1[24:0];
  assign operator_33_true_operator_33_true_or_tmp = (for_acc_1_tmp[6]) | operator_33_true_operator_33_true_and_tmp;
  assign nor_31_nl = ~(for_1_asn_sft_lpi_1_dfm_mx0 | (~ for_1_for_if_for_1_for_if_or_tmp));
  assign mux_nl = MUX_s_1_2_2(for_1_for_for_1_for_and_tmp, for_1_for_1_if_and_tmp,
      nor_31_nl);
  assign or_281_tmp = ((~ (mux_nl)) & for_1_for_1_and_1_tmp) | for_1_for_1_and_2_tmp;
  assign for_1_for_mux_5_nl = MUX_s_1_2_2(for_1_for_for_1_for_and_tmp, for_1_for_1_if_and_tmp,
      for_1_for_if_for_1_for_if_or_tmp);
  assign for_1_mux_1960_nl = MUX_s_1_2_2((for_1_for_mux_5_nl), for_1_for_for_1_for_and_tmp,
      for_1_asn_sft_lpi_1_dfm_mx0);
  assign for_1_and_1893_nl = (~ operator_33_true_operator_33_true_or_tmp) & for_1_or_tmp_1
      & (~ or_281_tmp);
  assign for_1_and_1894_nl = operator_33_true_operator_33_true_or_tmp & for_1_or_tmp_1
      & (~ or_281_tmp);
  assign and_32_nl = for_1_for_1_and_1_tmp & (~ or_281_tmp);
  assign for_1_mux1h_2098_tmp = MUX1HOT_v_2_4_2(2'b01, 2'b10, (signext_2_1(~ (for_1_mux_1960_nl))),
      lfst_exit_for_1_lpi_1_dfm_1, {(for_1_and_1893_nl) , (for_1_and_1894_nl) , (and_32_nl)
      , or_281_tmp});
  assign paramsIn_crt_lpi_1_dfm_12_0_mx0_12_11 = MUX_v_2_2_2((paramsIn_crt_lpi_1_dfm_12_0[12:11]),
      (paramsIn_rsci_idat_mxwt[12:11]), exitL_exit_for_1_sva);
  assign nl_for_acc_1_tmp = conv_u2s_6_7(for_i_6_0_lpi_1_dfm_1_5_0) + 7'b0000001;
  assign for_acc_1_tmp = nl_for_acc_1_tmp[6:0];
  assign operator_33_true_equal_tmp = (for_i_6_0_lpi_1_dfm_1_5_0) == (operator_11_false_2_acc_tmp[5:0]);
  assign operator_33_true_operator_33_true_and_tmp = operator_33_true_equal_tmp &
      (operator_11_false_2_acc_tmp[11:6]==6'b000000);
  assign for_1_mux_3_nl = MUX_v_11_2_2((paramsIn_crt_lpi_1_dfm_12_0[10:0]), (paramsIn_rsci_idat_mxwt[10:0]),
      exitL_exit_for_1_sva);
  assign nl_operator_11_false_2_acc_tmp = conv_u2s_11_12(for_1_mux_3_nl) + 12'b111111111111;
  assign operator_11_false_2_acc_tmp = nl_operator_11_false_2_acc_tmp[11:0];
  assign nand_7_nl = ~(main_stage_0_3 & for_1_and_1898_itm_1);
  assign for_1_mux_nl = MUX_v_25_2_2(tot_samples_in_img_mul_psp_sva_1, tot_samples_in_img_mul_psp_lpi_1,
      nand_7_nl);
  assign for_1_if_equal_tmp = (for_1_read_request_lpi_1[32:8]) == (for_1_mux_nl);
  assign for_1_for_1_if_and_tmp = (for_1_read_request_lpi_1[0]) & for_1_if_equal_tmp
      & (~((for_1_read_request_lpi_1[7:3]!=5'b00000))) & (~((for_1_read_request_lpi_1[36])
      | (for_1_read_request_lpi_1[35]) | (for_1_read_request_lpi_1[34]) | (for_1_read_request_lpi_1[33])
      | (for_1_read_request_lpi_1[2]) | (for_1_read_request_lpi_1[1]))) & (~((for_1_read_request_lpi_1[42:37]!=6'b000000)));
  assign for_1_not_3876_nl = ~ mux_89_cse;
  assign for_1_for_1_and_4_tmp = MUX_v_2_2_2(2'b00, for_1_mux1h_2098_tmp, (for_1_not_3876_nl));
  assign for_1_for_for_1_for_and_tmp = (~ operator_43_false_acc_itm_43) & exitL_exitL_exit_for_1_for_lpi_1;
  assign for_1_for_if_for_1_for_if_or_tmp = (operator_7_false_acc_tmp[6]) | ((~(for_1_for_if_unequal_tmp
      | (operator_11_false_2_acc_tmp[6]))) & (operator_11_false_2_acc_tmp[11:7]==5'b00000));
  assign nl_operator_7_false_acc_tmp = conv_u2u_6_7(for_1_for_quad_idx_lpi_1_dfm_5_0_1)
      + 7'b0000001;
  assign operator_7_false_acc_tmp = nl_operator_7_false_acc_tmp[6:0];
  assign for_1_for_1_for_nor_nl = ~(sfi_exit_for_1_lpi_1 | (~ for_1_for_for_1_for_and_1_tmp));
  assign for_1_for_quad_idx_lpi_1_dfm_5_0_1 = MUX_v_6_2_2(6'b000000, for_1_for_quad_idx_lpi_1_5_0,
      (for_1_for_1_for_nor_nl));
  assign for_1_for_if_unequal_tmp = for_1_for_quad_idx_lpi_1_dfm_5_0_1 != (operator_11_false_2_acc_tmp[5:0]);
  assign for_1_for_for_1_for_and_1_tmp = lfst_exitL_exit_for_1_for_lpi_1 & (~ exitL_exitL_exit_for_1_for_lpi_1);
  assign nl_operator_43_false_acc_nl = conv_u2s_43_44(for_1_read_request_lpi_1) +
      44'b11111111011111111111111111111111111111111111;
  assign operator_43_false_acc_nl = nl_operator_43_false_acc_nl[43:0];
  assign operator_43_false_acc_itm_43 = readslicef_44_1_43((operator_43_false_acc_nl));
  assign or_279_nl = (~ lfst_exitL_exit_for_1_for_lpi_1) | exitL_exitL_exit_for_1_for_lpi_1;
  assign for_1_asn_sft_lpi_1_dfm_mx0 = MUX_s_1_2_2(for_1_asn_sft_lpi_1, for_1_for_for_1_for_and_tmp,
      or_279_nl);
  assign for_1_for_1_and_1_tmp = (lfst_exit_for_1_lpi_1_dfm_1==2'b10);
  assign for_1_for_1_and_2_tmp = (lfst_exit_for_1_lpi_1_dfm_1==2'b11);
  assign paramsIn_crt_lpi_1_dfm_56_24_mx0 = MUX_v_33_2_2(paramsIn_crt_lpi_1_dfm_56_24,
      (paramsIn_rsci_idat_mxwt[45:13]), exitL_exit_for_1_sva);
  assign for_and_59_tmp = for_and_42_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_7_tmp = for_and_6_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_58_tmp = for_and_40_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_11_tmp = for_and_10_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_57_tmp = for_and_38_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_15_tmp = for_and_14_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_56_tmp = for_and_36_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_18_tmp = for_and_17_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_55_tmp = for_and_34_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_21_tmp = for_and_20_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_54_tmp = for_and_32_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_24_tmp = for_and_23_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_53_tmp = for_and_30_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_27_tmp = for_and_26_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_52_tmp = for_and_28_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_29_tmp = for_and_28_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_51_tmp = for_and_26_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_31_tmp = for_and_30_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_50_tmp = for_and_23_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_33_tmp = for_and_32_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_49_tmp = for_and_20_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_35_tmp = for_and_34_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_48_tmp = for_and_17_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_37_tmp = for_and_36_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_47_tmp = for_and_14_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_39_tmp = for_and_38_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_46_tmp = for_and_10_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_41_tmp = for_and_40_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_45_tmp = for_and_6_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_43_tmp = for_and_42_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[4]);
  assign for_and_44_tmp = for_and_2_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[4]));
  assign for_and_2_tmp = for_and_1_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_42_tmp = for_and_25_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_40_tmp = for_and_22_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_38_tmp = for_and_19_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_36_tmp = for_and_16_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_34_tmp = for_and_13_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_32_tmp = for_and_9_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_30_tmp = for_and_5_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_28_tmp = for_and_1_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[3]));
  assign for_and_26_tmp = for_and_25_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_23_tmp = for_and_22_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_20_tmp = for_and_19_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_17_tmp = for_and_16_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_14_tmp = for_and_13_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_10_tmp = for_and_9_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_6_tmp = for_and_5_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[3]);
  assign for_and_25_tmp = for_for_nor_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[2]));
  assign for_and_22_tmp = for_and_8_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[2]));
  assign for_and_19_tmp = for_and_4_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[2]));
  assign for_and_16_tmp = for_and_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[2]));
  assign for_and_13_tmp = for_for_nor_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[2]);
  assign for_and_9_tmp = for_and_8_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[2]);
  assign for_and_5_tmp = for_and_4_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[2]);
  assign for_and_1_tmp = for_and_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[2]);
  assign for_for_nor_tmp = ~((for_i_6_0_lpi_1_dfm_1_5_0[1:0]!=2'b00));
  assign for_and_8_tmp = (for_i_6_0_lpi_1_dfm_1_5_0[1:0]==2'b01);
  assign for_and_4_tmp = (for_i_6_0_lpi_1_dfm_1_5_0[1:0]==2'b10);
  assign for_and_tmp = (for_i_6_0_lpi_1_dfm_1_5_0[1:0]==2'b11);
  assign for_1_for_1_or_tmp = for_1_for_if_for_1_for_if_or_tmp | for_1_asn_sft_lpi_1_dfm_mx0;
  assign for_mux_nl = MUX_s_1_2_2(operator_33_true_operator_33_true_and_tmp, exit_for_sva,
      lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign for_1_for_1_nor_1894_nl = ~((for_mux_nl) | for_1_for_1_and_1_tmp | for_1_for_1_and_2_tmp);
  assign for_1_for_1_mux_76_tmp = MUX_v_6_2_2(for_i_6_0_lpi_1_dfm_1_5_0, (for_acc_1_tmp[5:0]),
      for_1_for_1_nor_1894_nl);
  assign and_dcpl_6 = (operator_11_false_2_acc_tmp[11:6]==6'b000000) & operator_33_true_equal_tmp;
  assign and_dcpl_7 = (and_dcpl_6 | (for_acc_1_tmp[6])) & (~ (lfst_exit_for_1_lpi_1_dfm_1[1]))
      & main_stage_0_2;
  assign or_tmp_5 = exitL_exitL_exit_for_1_for_lpi_1 | for_1_or_tmp_1 | sfi_exit_for_1_lpi_1
      | (~ lfst_exitL_exit_for_1_for_lpi_1) | for_1_asn_sft_lpi_1;
  assign nor_tmp_2 = lfst_exitL_exit_for_1_for_lpi_1 & for_1_asn_sft_lpi_1;
  assign or_8_nl = for_1_or_tmp_1 | nor_tmp_2;
  assign or_7_nl = (~ operator_43_false_acc_itm_43) | for_1_or_tmp_1;
  assign mux_tmp_2 = MUX_s_1_2_2((or_8_nl), (or_7_nl), exitL_exitL_exit_for_1_for_lpi_1);
  assign or_19_nl = (((for_1_for_1_mux_76_tmp!=6'b000000)) & (for_1_mux1h_2098_tmp[0]))
      | (for_1_mux1h_2098_tmp[1]);
  assign mux_tmp_9 = MUX_s_1_2_2((~ exitL_exit_for_1_sva), (or_19_nl), main_stage_0_2);
  assign or_22_nl = (for_1_for_1_mux_76_tmp!=6'b000001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_10 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_22_nl), main_stage_0_2);
  assign or_24_nl = (for_1_for_1_mux_76_tmp!=6'b000010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_11 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_24_nl), main_stage_0_2);
  assign or_26_nl = (for_1_for_1_mux_76_tmp!=6'b000011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_12 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_26_nl), main_stage_0_2);
  assign or_28_nl = (for_1_for_1_mux_76_tmp!=6'b000100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_13 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_28_nl), main_stage_0_2);
  assign or_30_nl = (for_1_for_1_mux_76_tmp!=6'b000101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_14 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_30_nl), main_stage_0_2);
  assign or_32_nl = (for_1_for_1_mux_76_tmp!=6'b000110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_15 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_32_nl), main_stage_0_2);
  assign or_34_nl = (for_1_for_1_mux_76_tmp!=6'b000111) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_16 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_34_nl), main_stage_0_2);
  assign or_36_nl = (for_1_for_1_mux_76_tmp!=6'b001000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_17 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_36_nl), main_stage_0_2);
  assign or_38_nl = (for_1_for_1_mux_76_tmp!=6'b001001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_18 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_38_nl), main_stage_0_2);
  assign or_40_nl = (for_1_for_1_mux_76_tmp!=6'b001010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_19 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_40_nl), main_stage_0_2);
  assign or_42_nl = (for_1_for_1_mux_76_tmp!=6'b001011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_20 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_42_nl), main_stage_0_2);
  assign or_44_nl = (for_1_for_1_mux_76_tmp!=6'b001100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_21 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_44_nl), main_stage_0_2);
  assign or_46_nl = (for_1_for_1_mux_76_tmp!=6'b001101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_22 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_46_nl), main_stage_0_2);
  assign or_48_nl = (for_1_for_1_mux_76_tmp!=6'b001110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_23 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_48_nl), main_stage_0_2);
  assign or_50_nl = (for_1_for_1_mux_76_tmp!=6'b001111) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_24 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_50_nl), main_stage_0_2);
  assign or_52_nl = (for_1_for_1_mux_76_tmp!=6'b010000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_25 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_52_nl), main_stage_0_2);
  assign or_54_nl = (for_1_for_1_mux_76_tmp!=6'b010001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_26 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_54_nl), main_stage_0_2);
  assign or_56_nl = (for_1_for_1_mux_76_tmp!=6'b010010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_27 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_56_nl), main_stage_0_2);
  assign or_58_nl = (for_1_for_1_mux_76_tmp!=6'b010011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_28 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_58_nl), main_stage_0_2);
  assign or_60_nl = (for_1_for_1_mux_76_tmp!=6'b010100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_29 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_60_nl), main_stage_0_2);
  assign or_62_nl = (for_1_for_1_mux_76_tmp!=6'b010101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_30 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_62_nl), main_stage_0_2);
  assign or_64_nl = (for_1_for_1_mux_76_tmp!=6'b010110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_31 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_64_nl), main_stage_0_2);
  assign or_66_nl = (for_1_for_1_mux_76_tmp!=6'b010111) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_32 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_66_nl), main_stage_0_2);
  assign or_68_nl = (for_1_for_1_mux_76_tmp!=6'b011000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_33 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_68_nl), main_stage_0_2);
  assign or_70_nl = (for_1_for_1_mux_76_tmp!=6'b011001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_34 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_70_nl), main_stage_0_2);
  assign or_72_nl = (for_1_for_1_mux_76_tmp!=6'b011010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_35 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_72_nl), main_stage_0_2);
  assign or_74_nl = (for_1_for_1_mux_76_tmp!=6'b011011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_36 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_74_nl), main_stage_0_2);
  assign or_76_nl = (for_1_for_1_mux_76_tmp!=6'b011100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_37 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_76_nl), main_stage_0_2);
  assign or_78_nl = (for_1_for_1_mux_76_tmp!=6'b011101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_38 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_78_nl), main_stage_0_2);
  assign or_80_nl = (for_1_for_1_mux_76_tmp!=6'b011110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_39 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_80_nl), main_stage_0_2);
  assign nand_1_nl = ~((for_1_for_1_mux_76_tmp==6'b011111) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_40 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_1_nl), main_stage_0_2);
  assign or_84_nl = (for_1_for_1_mux_76_tmp!=6'b100000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_41 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_84_nl), main_stage_0_2);
  assign or_86_nl = (for_1_for_1_mux_76_tmp!=6'b100001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_42 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_86_nl), main_stage_0_2);
  assign or_88_nl = (for_1_for_1_mux_76_tmp!=6'b100010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_43 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_88_nl), main_stage_0_2);
  assign or_90_nl = (for_1_for_1_mux_76_tmp!=6'b100011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_44 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_90_nl), main_stage_0_2);
  assign or_92_nl = (for_1_for_1_mux_76_tmp!=6'b100100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_45 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_92_nl), main_stage_0_2);
  assign or_94_nl = (for_1_for_1_mux_76_tmp!=6'b100101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_46 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_94_nl), main_stage_0_2);
  assign or_96_nl = (for_1_for_1_mux_76_tmp!=6'b100110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_47 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_96_nl), main_stage_0_2);
  assign or_98_nl = (for_1_for_1_mux_76_tmp!=6'b100111) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_48 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_98_nl), main_stage_0_2);
  assign or_100_nl = (for_1_for_1_mux_76_tmp!=6'b101000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_49 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_100_nl), main_stage_0_2);
  assign or_102_nl = (for_1_for_1_mux_76_tmp!=6'b101001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_50 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_102_nl), main_stage_0_2);
  assign or_104_nl = (for_1_for_1_mux_76_tmp!=6'b101010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_51 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_104_nl), main_stage_0_2);
  assign or_106_nl = (for_1_for_1_mux_76_tmp!=6'b101011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_52 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_106_nl), main_stage_0_2);
  assign or_108_nl = (for_1_for_1_mux_76_tmp!=6'b101100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_53 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_108_nl), main_stage_0_2);
  assign or_110_nl = (for_1_for_1_mux_76_tmp!=6'b101101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_54 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_110_nl), main_stage_0_2);
  assign or_112_nl = (for_1_for_1_mux_76_tmp!=6'b101110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_55 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_112_nl), main_stage_0_2);
  assign nand_2_nl = ~((for_1_for_1_mux_76_tmp==6'b101111) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_56 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_2_nl), main_stage_0_2);
  assign or_116_nl = (for_1_for_1_mux_76_tmp!=6'b110000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_57 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_116_nl), main_stage_0_2);
  assign or_118_nl = (for_1_for_1_mux_76_tmp!=6'b110001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_58 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_118_nl), main_stage_0_2);
  assign or_120_nl = (for_1_for_1_mux_76_tmp!=6'b110010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_59 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_120_nl), main_stage_0_2);
  assign or_122_nl = (for_1_for_1_mux_76_tmp!=6'b110011) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_60 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_122_nl), main_stage_0_2);
  assign or_124_nl = (for_1_for_1_mux_76_tmp!=6'b110100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_61 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_124_nl), main_stage_0_2);
  assign or_126_nl = (for_1_for_1_mux_76_tmp!=6'b110101) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_62 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_126_nl), main_stage_0_2);
  assign or_128_nl = (for_1_for_1_mux_76_tmp!=6'b110110) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_63 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_128_nl), main_stage_0_2);
  assign nand_3_nl = ~((for_1_for_1_mux_76_tmp==6'b110111) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_64 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_3_nl), main_stage_0_2);
  assign or_132_nl = (for_1_for_1_mux_76_tmp!=6'b111000) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_65 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_132_nl), main_stage_0_2);
  assign or_134_nl = (for_1_for_1_mux_76_tmp!=6'b111001) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_66 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_134_nl), main_stage_0_2);
  assign or_136_nl = (for_1_for_1_mux_76_tmp!=6'b111010) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_67 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_136_nl), main_stage_0_2);
  assign nand_4_nl = ~((for_1_for_1_mux_76_tmp==6'b111011) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_68 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_4_nl), main_stage_0_2);
  assign or_140_nl = (for_1_for_1_mux_76_tmp!=6'b111100) | (for_1_mux1h_2098_tmp!=2'b01);
  assign mux_tmp_69 = MUX_s_1_2_2(exitL_exit_for_1_sva, (or_140_nl), main_stage_0_2);
  assign nand_5_nl = ~((for_1_for_1_mux_76_tmp==6'b111101) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_70 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_5_nl), main_stage_0_2);
  assign nand_6_nl = ~((for_1_for_1_mux_76_tmp==6'b111110) & (for_1_mux1h_2098_tmp==2'b01));
  assign mux_tmp_71 = MUX_s_1_2_2(exitL_exit_for_1_sva, (nand_6_nl), main_stage_0_2);
  assign or_tmp_161 = for_1_for_if_unequal_tmp | (operator_11_false_2_acc_tmp[11:6]!=6'b000000);
  assign or_tmp_162 = nor_tmp_2 | (~ or_tmp_161);
  assign or_dcpl_2 = (lfst_exit_for_1_lpi_1_dfm_1[1]) | (~ main_stage_0_2);
  assign or_dcpl_12 = (lfst_exit_for_1_lpi_1_dfm_1!=2'b10) | (~ main_stage_0_2);
  assign mux_88_nl = MUX_s_1_2_2(nor_tmp_2, (~ operator_43_false_acc_itm_43), exitL_exitL_exit_for_1_for_lpi_1);
  assign or_dcpl_13 = (mux_88_nl) | or_dcpl_12;
  assign or_dcpl_14 = (for_i_6_0_lpi_1_dfm_1_5_0[5:4]!=2'b00);
  assign or_dcpl_15 = (for_i_6_0_lpi_1_dfm_1_5_0[3:2]!=2'b00);
  assign or_dcpl_16 = or_dcpl_15 | or_dcpl_14;
  assign or_dcpl_18 = or_dcpl_2 | (for_i_6_0_lpi_1_dfm_1_5_0[1:0]!=2'b00);
  assign or_dcpl_21 = or_dcpl_2 | (for_i_6_0_lpi_1_dfm_1_5_0[1:0]!=2'b01);
  assign or_dcpl_24 = or_dcpl_2 | (for_i_6_0_lpi_1_dfm_1_5_0[1:0]!=2'b10);
  assign or_dcpl_27 = or_dcpl_2 | (for_i_6_0_lpi_1_dfm_1_5_0[1:0]!=2'b11);
  assign or_dcpl_29 = (for_i_6_0_lpi_1_dfm_1_5_0[3:2]!=2'b01);
  assign or_dcpl_30 = or_dcpl_29 | or_dcpl_14;
  assign or_dcpl_35 = (for_i_6_0_lpi_1_dfm_1_5_0[3:2]!=2'b10);
  assign or_dcpl_36 = or_dcpl_35 | or_dcpl_14;
  assign or_dcpl_41 = ~((for_i_6_0_lpi_1_dfm_1_5_0[3:2]==2'b11));
  assign or_dcpl_42 = or_dcpl_41 | or_dcpl_14;
  assign or_dcpl_47 = (for_i_6_0_lpi_1_dfm_1_5_0[5:4]!=2'b01);
  assign or_dcpl_48 = or_dcpl_15 | or_dcpl_47;
  assign or_dcpl_53 = or_dcpl_29 | or_dcpl_47;
  assign or_dcpl_58 = or_dcpl_35 | or_dcpl_47;
  assign or_dcpl_63 = or_dcpl_41 | or_dcpl_47;
  assign or_dcpl_68 = (for_i_6_0_lpi_1_dfm_1_5_0[5:4]!=2'b10);
  assign or_dcpl_69 = or_dcpl_15 | or_dcpl_68;
  assign or_dcpl_74 = or_dcpl_29 | or_dcpl_68;
  assign or_dcpl_79 = or_dcpl_35 | or_dcpl_68;
  assign or_dcpl_84 = or_dcpl_41 | or_dcpl_68;
  assign or_dcpl_89 = ~((for_i_6_0_lpi_1_dfm_1_5_0[5:4]==2'b11));
  assign or_dcpl_90 = or_dcpl_15 | or_dcpl_89;
  assign or_dcpl_95 = or_dcpl_29 | or_dcpl_89;
  assign or_dcpl_100 = or_dcpl_35 | or_dcpl_89;
  assign or_dcpl_105 = or_dcpl_41 | or_dcpl_89;
  assign mux_tmp_89 = MUX_s_1_2_2((~ exitL_exit_for_1_sva), or_1_cse, main_stage_0_2);
  assign or_287_nl = (operator_11_false_2_acc_tmp[11:6]!=6'b000000) | for_1_for_if_unequal_tmp
      | (~ (for_1_read_request_lpi_1[0])) | (~ for_1_if_equal_tmp) | (for_1_read_request_lpi_1[7])
      | (for_1_read_request_lpi_1[6]) | (for_1_read_request_lpi_1[5]) | (for_1_read_request_lpi_1[4])
      | (for_1_read_request_lpi_1[3]) | (for_1_read_request_lpi_1[36]) | (for_1_read_request_lpi_1[35])
      | (for_1_read_request_lpi_1[34]) | (for_1_read_request_lpi_1[33]) | (for_1_read_request_lpi_1[2])
      | (for_1_read_request_lpi_1[1]) | (for_1_read_request_lpi_1[42]) | (for_1_read_request_lpi_1[41])
      | (for_1_read_request_lpi_1[40]) | (for_1_read_request_lpi_1[39]) | (for_1_read_request_lpi_1[38])
      | (for_1_read_request_lpi_1[37]);
  assign or_286_nl = (~ (for_1_read_request_lpi_1[0])) | (~ for_1_if_equal_tmp) |
      (for_1_read_request_lpi_1[7]) | (for_1_read_request_lpi_1[6]) | (for_1_read_request_lpi_1[5])
      | (for_1_read_request_lpi_1[4]) | (for_1_read_request_lpi_1[3]) | (for_1_read_request_lpi_1[36])
      | (for_1_read_request_lpi_1[35]) | (for_1_read_request_lpi_1[34]) | (for_1_read_request_lpi_1[33])
      | (for_1_read_request_lpi_1[2]) | (for_1_read_request_lpi_1[1]) | (for_1_read_request_lpi_1[42])
      | (for_1_read_request_lpi_1[41]) | (for_1_read_request_lpi_1[40]) | (for_1_read_request_lpi_1[39])
      | (for_1_read_request_lpi_1[38]) | (for_1_read_request_lpi_1[37]);
  assign mux_tmp_91 = MUX_s_1_2_2((or_287_nl), (or_286_nl), operator_7_false_acc_tmp[6]);
  assign or_288_nl = nor_tmp_2 | mux_tmp_91;
  assign and_38_nl = operator_43_false_acc_itm_43 & mux_tmp_91;
  assign mux_95_nl = MUX_s_1_2_2((or_288_nl), (and_38_nl), exitL_exitL_exit_for_1_for_lpi_1);
  assign or_289_nl = (lfst_exit_for_1_lpi_1_dfm_1[0]) | (mux_95_nl);
  assign mux_tmp_93 = MUX_s_1_2_2((~ for_1_or_tmp_1), (or_289_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign or_302_cse = (~ (lfst_exit_for_1_lpi_1_dfm_1[1])) | for_1_or_tmp_1;
  assign nor_tmp_14 = or_302_cse & (for_acc_1_tmp[6]);
  assign or_tmp_183 = operator_33_true_equal_tmp | (for_acc_1_tmp[6]);
  assign and_tmp_2 = or_302_cse & or_tmp_183;
  assign nor_tmp_15 = for_1_or_tmp_1 & (for_acc_1_tmp[6]);
  assign and_tmp_3 = for_1_or_tmp_1 & or_tmp_183;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      tot_samples_in_img_mul_psp_lpi_1 <= 25'b0000000000000000000000000;
    end
    else if ( run_wen & ((((~((~((operator_11_false_2_acc_tmp[11:6]!=6'b000000) |
        (~ operator_33_true_equal_tmp))) | (for_acc_1_tmp[6]))) | or_dcpl_2) & main_stage_0_3
        & for_1_and_1898_itm_1) | and_dcpl_7) ) begin
      tot_samples_in_img_mul_psp_lpi_1 <= MUX_v_25_2_2(tot_samples_in_img_mul_psp_sva_1,
          ({3'b000 , (pixels_in_img_mul_nl)}), and_dcpl_7);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_2_false_2_operator_2_false_2_and_mdf_sva_1 <= 1'b0;
      operator_2_false_1_operator_2_false_1_and_mdf_sva_1 <= 1'b0;
      operator_2_false_operator_2_false_nor_mdf_sva_1 <= 1'b0;
    end
    else if ( qelse_qelse_and_cse ) begin
      operator_2_false_2_operator_2_false_2_and_mdf_sva_1 <= (paramsIn_crt_lpi_1_dfm_12_0_mx0_12_11==2'b10);
      operator_2_false_1_operator_2_false_1_and_mdf_sva_1 <= (paramsIn_crt_lpi_1_dfm_12_0_mx0_12_11==2'b01);
      operator_2_false_operator_2_false_nor_mdf_sva_1 <= ~((paramsIn_crt_lpi_1_dfm_12_0_mx0_12_11!=2'b00));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_1_and_1898_itm_1 <= 1'b0;
      reg_quads_out_rsci_oswt_cse <= 1'b0;
      reg_paramsIn_rsci_oswt_cse <= 1'b0;
      reg_quads_in_rsci_oswt_cse <= 1'b0;
      for_1_or_tmp_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
    end
    else if ( run_wen ) begin
      for_1_and_1898_itm_1 <= operator_33_true_operator_33_true_or_tmp & (~(for_1_for_1_and_1_tmp
          | for_1_for_1_and_2_tmp));
      reg_quads_out_rsci_oswt_cse <= ~ or_dcpl_13;
      reg_paramsIn_rsci_oswt_cse <= mux_89_cse;
      reg_quads_in_rsci_oswt_cse <= MUX_s_1_2_2(exitL_exit_for_1_sva, (~ (for_1_mux1h_2098_tmp[1])),
          main_stage_0_2);
      for_1_or_tmp_1 <= ((for_1_for_1_and_4_tmp==2'b01)) | (~((for_1_for_1_and_4_tmp!=2'b00)));
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_out_rsci_idat_376_352 <= 25'b0000000000000000000000000;
      quads_out_rsci_idat_11_0 <= 12'b000000000000;
      quads_out_rsci_idat_351_350 <= 2'b00;
      quads_out_rsci_idat_23_12 <= 12'b000000000000;
      quads_out_rsci_idat_349_323 <= 27'b000000000000000000000000000;
      quads_out_rsci_idat_31_24 <= 8'b00000000;
      quads_out_rsci_idat_322_320 <= 3'b000;
      quads_out_rsci_idat_35_32 <= 4'b0000;
      quads_out_rsci_idat_319_296 <= 24'b000000000000000000000000;
      quads_out_rsci_idat_47_36 <= 12'b000000000000;
      quads_out_rsci_idat_295_288 <= 8'b00000000;
      quads_out_rsci_idat_59_48 <= 12'b000000000000;
      quads_out_rsci_idat_287_265 <= 23'b00000000000000000000000;
      quads_out_rsci_idat_63_60 <= 4'b0000;
      quads_out_rsci_idat_264_256 <= 9'b000000000;
      quads_out_rsci_idat_71_64 <= 8'b00000000;
      quads_out_rsci_idat_255_240 <= 16'b0000000000000000;
      quads_out_rsci_idat_83_72 <= 12'b000000000000;
      quads_out_rsci_idat_239_224 <= 16'b0000000000000000;
      quads_out_rsci_idat_95_84 <= 12'b000000000000;
      quads_out_rsci_idat_223_215 <= 9'b000000000;
      quads_out_rsci_idat_107_96 <= 12'b000000000000;
      quads_out_rsci_idat_214_192 <= 23'b00000000000000000000000;
      quads_out_rsci_idat_110_108 <= 3'b000;
      quads_out_rsci_idat_191_190 <= 2'b00;
      quads_out_rsci_idat_111 <= 1'b0;
      quads_out_rsci_idat_189_164 <= 26'b00000000000000000000000000;
      quads_out_rsci_idat_127_112 <= 16'b0000000000000000;
      quads_out_rsci_idat_163_160 <= 4'b0000;
      quads_out_rsci_idat_137_128 <= 10'b0000000000;
      quads_out_rsci_idat_159_138 <= 22'b0000000000000000000000;
    end
    else if ( quads_out_and_cse ) begin
      quads_out_rsci_idat_376_352 <= MUX_v_25_64_2(buffer_bank11_data_0_lpi_1, buffer_bank11_data_1_lpi_1,
          buffer_bank11_data_2_lpi_1, buffer_bank11_data_3_lpi_1, buffer_bank11_data_4_lpi_1,
          buffer_bank11_data_5_lpi_1, buffer_bank11_data_6_lpi_1, buffer_bank11_data_7_lpi_1,
          buffer_bank11_data_8_lpi_1, buffer_bank11_data_9_lpi_1, buffer_bank11_data_10_lpi_1,
          buffer_bank11_data_11_lpi_1, buffer_bank11_data_12_lpi_1, buffer_bank11_data_13_lpi_1,
          buffer_bank11_data_14_lpi_1, buffer_bank11_data_15_lpi_1, buffer_bank11_data_16_lpi_1,
          buffer_bank11_data_17_lpi_1, buffer_bank11_data_18_lpi_1, buffer_bank11_data_19_lpi_1,
          buffer_bank11_data_20_lpi_1, buffer_bank11_data_21_lpi_1, buffer_bank11_data_22_lpi_1,
          buffer_bank11_data_23_lpi_1, buffer_bank11_data_24_lpi_1, buffer_bank11_data_25_lpi_1,
          buffer_bank11_data_26_lpi_1, buffer_bank11_data_27_lpi_1, buffer_bank11_data_28_lpi_1,
          buffer_bank11_data_29_lpi_1, buffer_bank11_data_30_lpi_1, buffer_bank11_data_31_lpi_1,
          buffer_bank11_data_32_lpi_1, buffer_bank11_data_33_lpi_1, buffer_bank11_data_34_lpi_1,
          buffer_bank11_data_35_lpi_1, buffer_bank11_data_36_lpi_1, buffer_bank11_data_37_lpi_1,
          buffer_bank11_data_38_lpi_1, buffer_bank11_data_39_lpi_1, buffer_bank11_data_40_lpi_1,
          buffer_bank11_data_41_lpi_1, buffer_bank11_data_42_lpi_1, buffer_bank11_data_43_lpi_1,
          buffer_bank11_data_44_lpi_1, buffer_bank11_data_45_lpi_1, buffer_bank11_data_46_lpi_1,
          buffer_bank11_data_47_lpi_1, buffer_bank11_data_48_lpi_1, buffer_bank11_data_49_lpi_1,
          buffer_bank11_data_50_lpi_1, buffer_bank11_data_51_lpi_1, buffer_bank11_data_52_lpi_1,
          buffer_bank11_data_53_lpi_1, buffer_bank11_data_54_lpi_1, buffer_bank11_data_55_lpi_1,
          buffer_bank11_data_56_lpi_1, buffer_bank11_data_57_lpi_1, buffer_bank11_data_58_lpi_1,
          buffer_bank11_data_59_lpi_1, buffer_bank11_data_60_lpi_1, buffer_bank11_data_61_lpi_1,
          buffer_bank11_data_62_lpi_1, (quads_in_crt_lpi_1[376:352]), for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_11_0 <= MUX_v_12_64_2(buffer_bank0_data_0_11_0_lpi_1, buffer_bank0_data_1_11_0_lpi_1,
          buffer_bank0_data_2_11_0_lpi_1, buffer_bank0_data_3_11_0_lpi_1, buffer_bank0_data_4_11_0_lpi_1,
          buffer_bank0_data_5_11_0_lpi_1, buffer_bank0_data_6_11_0_lpi_1, buffer_bank0_data_7_11_0_lpi_1,
          buffer_bank0_data_8_11_0_lpi_1, buffer_bank0_data_9_11_0_lpi_1, buffer_bank0_data_10_11_0_lpi_1,
          buffer_bank0_data_11_11_0_lpi_1, buffer_bank0_data_12_11_0_lpi_1, buffer_bank0_data_13_11_0_lpi_1,
          buffer_bank0_data_14_11_0_lpi_1, buffer_bank0_data_15_11_0_lpi_1, buffer_bank0_data_16_11_0_lpi_1,
          buffer_bank0_data_17_11_0_lpi_1, buffer_bank0_data_18_11_0_lpi_1, buffer_bank0_data_19_11_0_lpi_1,
          buffer_bank0_data_20_11_0_lpi_1, buffer_bank0_data_21_11_0_lpi_1, buffer_bank0_data_22_11_0_lpi_1,
          buffer_bank0_data_23_11_0_lpi_1, buffer_bank0_data_24_11_0_lpi_1, buffer_bank0_data_25_11_0_lpi_1,
          buffer_bank0_data_26_11_0_lpi_1, buffer_bank0_data_27_11_0_lpi_1, buffer_bank0_data_28_11_0_lpi_1,
          buffer_bank0_data_29_11_0_lpi_1, buffer_bank0_data_30_11_0_lpi_1, buffer_bank0_data_31_11_0_lpi_1,
          buffer_bank0_data_32_11_0_lpi_1, buffer_bank0_data_33_11_0_lpi_1, buffer_bank0_data_34_11_0_lpi_1,
          buffer_bank0_data_35_11_0_lpi_1, buffer_bank0_data_36_11_0_lpi_1, buffer_bank0_data_37_11_0_lpi_1,
          buffer_bank0_data_38_11_0_lpi_1, buffer_bank0_data_39_11_0_lpi_1, buffer_bank0_data_40_11_0_lpi_1,
          buffer_bank0_data_41_11_0_lpi_1, buffer_bank0_data_42_11_0_lpi_1, buffer_bank0_data_43_11_0_lpi_1,
          buffer_bank0_data_44_11_0_lpi_1, buffer_bank0_data_45_11_0_lpi_1, buffer_bank0_data_46_11_0_lpi_1,
          buffer_bank0_data_47_11_0_lpi_1, buffer_bank0_data_48_11_0_lpi_1, buffer_bank0_data_49_11_0_lpi_1,
          buffer_bank0_data_50_11_0_lpi_1, buffer_bank0_data_51_11_0_lpi_1, buffer_bank0_data_52_11_0_lpi_1,
          buffer_bank0_data_53_11_0_lpi_1, buffer_bank0_data_54_11_0_lpi_1, buffer_bank0_data_55_11_0_lpi_1,
          buffer_bank0_data_56_11_0_lpi_1, buffer_bank0_data_57_11_0_lpi_1, buffer_bank0_data_58_11_0_lpi_1,
          buffer_bank0_data_59_11_0_lpi_1, buffer_bank0_data_60_11_0_lpi_1, buffer_bank0_data_61_11_0_lpi_1,
          buffer_bank0_data_62_11_0_lpi_1, (quads_in_crt_lpi_1[11:0]), for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_351_350 <= MUX_v_2_64_2(buffer_bank10_data_0_31_30_lpi_1,
          buffer_bank10_data_1_31_30_lpi_1, buffer_bank10_data_2_31_30_lpi_1, buffer_bank10_data_3_31_30_lpi_1,
          buffer_bank10_data_4_31_30_lpi_1, buffer_bank10_data_5_31_30_lpi_1, buffer_bank10_data_6_31_30_lpi_1,
          buffer_bank10_data_7_31_30_lpi_1, buffer_bank10_data_8_31_30_lpi_1, buffer_bank10_data_9_31_30_lpi_1,
          buffer_bank10_data_10_31_30_lpi_1, buffer_bank10_data_11_31_30_lpi_1, buffer_bank10_data_12_31_30_lpi_1,
          buffer_bank10_data_13_31_30_lpi_1, buffer_bank10_data_14_31_30_lpi_1, buffer_bank10_data_15_31_30_lpi_1,
          buffer_bank10_data_16_31_30_lpi_1, buffer_bank10_data_17_31_30_lpi_1, buffer_bank10_data_18_31_30_lpi_1,
          buffer_bank10_data_19_31_30_lpi_1, buffer_bank10_data_20_31_30_lpi_1, buffer_bank10_data_21_31_30_lpi_1,
          buffer_bank10_data_22_31_30_lpi_1, buffer_bank10_data_23_31_30_lpi_1, buffer_bank10_data_24_31_30_lpi_1,
          buffer_bank10_data_25_31_30_lpi_1, buffer_bank10_data_26_31_30_lpi_1, buffer_bank10_data_27_31_30_lpi_1,
          buffer_bank10_data_28_31_30_lpi_1, buffer_bank10_data_29_31_30_lpi_1, buffer_bank10_data_30_31_30_lpi_1,
          buffer_bank10_data_31_31_30_lpi_1, buffer_bank10_data_32_31_30_lpi_1, buffer_bank10_data_33_31_30_lpi_1,
          buffer_bank10_data_34_31_30_lpi_1, buffer_bank10_data_35_31_30_lpi_1, buffer_bank10_data_36_31_30_lpi_1,
          buffer_bank10_data_37_31_30_lpi_1, buffer_bank10_data_38_31_30_lpi_1, buffer_bank10_data_39_31_30_lpi_1,
          buffer_bank10_data_40_31_30_lpi_1, buffer_bank10_data_41_31_30_lpi_1, buffer_bank10_data_42_31_30_lpi_1,
          buffer_bank10_data_43_31_30_lpi_1, buffer_bank10_data_44_31_30_lpi_1, buffer_bank10_data_45_31_30_lpi_1,
          buffer_bank10_data_46_31_30_lpi_1, buffer_bank10_data_47_31_30_lpi_1, buffer_bank10_data_48_31_30_lpi_1,
          buffer_bank10_data_49_31_30_lpi_1, buffer_bank10_data_50_31_30_lpi_1, buffer_bank10_data_51_31_30_lpi_1,
          buffer_bank10_data_52_31_30_lpi_1, buffer_bank10_data_53_31_30_lpi_1, buffer_bank10_data_54_31_30_lpi_1,
          buffer_bank10_data_55_31_30_lpi_1, buffer_bank10_data_56_31_30_lpi_1, buffer_bank10_data_57_31_30_lpi_1,
          buffer_bank10_data_58_31_30_lpi_1, buffer_bank10_data_59_31_30_lpi_1, buffer_bank10_data_60_31_30_lpi_1,
          buffer_bank10_data_61_31_30_lpi_1, buffer_bank10_data_62_31_30_lpi_1, (quads_in_crt_lpi_1[351:350]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_23_12 <= MUX_v_12_64_2(buffer_bank0_data_0_23_12_lpi_1,
          buffer_bank0_data_1_23_12_lpi_1, buffer_bank0_data_2_23_12_lpi_1, buffer_bank0_data_3_23_12_lpi_1,
          buffer_bank0_data_4_23_12_lpi_1, buffer_bank0_data_5_23_12_lpi_1, buffer_bank0_data_6_23_12_lpi_1,
          buffer_bank0_data_7_23_12_lpi_1, buffer_bank0_data_8_23_12_lpi_1, buffer_bank0_data_9_23_12_lpi_1,
          buffer_bank0_data_10_23_12_lpi_1, buffer_bank0_data_11_23_12_lpi_1, buffer_bank0_data_12_23_12_lpi_1,
          buffer_bank0_data_13_23_12_lpi_1, buffer_bank0_data_14_23_12_lpi_1, buffer_bank0_data_15_23_12_lpi_1,
          buffer_bank0_data_16_23_12_lpi_1, buffer_bank0_data_17_23_12_lpi_1, buffer_bank0_data_18_23_12_lpi_1,
          buffer_bank0_data_19_23_12_lpi_1, buffer_bank0_data_20_23_12_lpi_1, buffer_bank0_data_21_23_12_lpi_1,
          buffer_bank0_data_22_23_12_lpi_1, buffer_bank0_data_23_23_12_lpi_1, buffer_bank0_data_24_23_12_lpi_1,
          buffer_bank0_data_25_23_12_lpi_1, buffer_bank0_data_26_23_12_lpi_1, buffer_bank0_data_27_23_12_lpi_1,
          buffer_bank0_data_28_23_12_lpi_1, buffer_bank0_data_29_23_12_lpi_1, buffer_bank0_data_30_23_12_lpi_1,
          buffer_bank0_data_31_23_12_lpi_1, buffer_bank0_data_32_23_12_lpi_1, buffer_bank0_data_33_23_12_lpi_1,
          buffer_bank0_data_34_23_12_lpi_1, buffer_bank0_data_35_23_12_lpi_1, buffer_bank0_data_36_23_12_lpi_1,
          buffer_bank0_data_37_23_12_lpi_1, buffer_bank0_data_38_23_12_lpi_1, buffer_bank0_data_39_23_12_lpi_1,
          buffer_bank0_data_40_23_12_lpi_1, buffer_bank0_data_41_23_12_lpi_1, buffer_bank0_data_42_23_12_lpi_1,
          buffer_bank0_data_43_23_12_lpi_1, buffer_bank0_data_44_23_12_lpi_1, buffer_bank0_data_45_23_12_lpi_1,
          buffer_bank0_data_46_23_12_lpi_1, buffer_bank0_data_47_23_12_lpi_1, buffer_bank0_data_48_23_12_lpi_1,
          buffer_bank0_data_49_23_12_lpi_1, buffer_bank0_data_50_23_12_lpi_1, buffer_bank0_data_51_23_12_lpi_1,
          buffer_bank0_data_52_23_12_lpi_1, buffer_bank0_data_53_23_12_lpi_1, buffer_bank0_data_54_23_12_lpi_1,
          buffer_bank0_data_55_23_12_lpi_1, buffer_bank0_data_56_23_12_lpi_1, buffer_bank0_data_57_23_12_lpi_1,
          buffer_bank0_data_58_23_12_lpi_1, buffer_bank0_data_59_23_12_lpi_1, buffer_bank0_data_60_23_12_lpi_1,
          buffer_bank0_data_61_23_12_lpi_1, buffer_bank0_data_62_23_12_lpi_1, (quads_in_crt_lpi_1[23:12]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_349_323 <= MUX_v_27_64_2(buffer_bank10_data_0_29_3_lpi_1,
          buffer_bank10_data_1_29_3_lpi_1, buffer_bank10_data_2_29_3_lpi_1, buffer_bank10_data_3_29_3_lpi_1,
          buffer_bank10_data_4_29_3_lpi_1, buffer_bank10_data_5_29_3_lpi_1, buffer_bank10_data_6_29_3_lpi_1,
          buffer_bank10_data_7_29_3_lpi_1, buffer_bank10_data_8_29_3_lpi_1, buffer_bank10_data_9_29_3_lpi_1,
          buffer_bank10_data_10_29_3_lpi_1, buffer_bank10_data_11_29_3_lpi_1, buffer_bank10_data_12_29_3_lpi_1,
          buffer_bank10_data_13_29_3_lpi_1, buffer_bank10_data_14_29_3_lpi_1, buffer_bank10_data_15_29_3_lpi_1,
          buffer_bank10_data_16_29_3_lpi_1, buffer_bank10_data_17_29_3_lpi_1, buffer_bank10_data_18_29_3_lpi_1,
          buffer_bank10_data_19_29_3_lpi_1, buffer_bank10_data_20_29_3_lpi_1, buffer_bank10_data_21_29_3_lpi_1,
          buffer_bank10_data_22_29_3_lpi_1, buffer_bank10_data_23_29_3_lpi_1, buffer_bank10_data_24_29_3_lpi_1,
          buffer_bank10_data_25_29_3_lpi_1, buffer_bank10_data_26_29_3_lpi_1, buffer_bank10_data_27_29_3_lpi_1,
          buffer_bank10_data_28_29_3_lpi_1, buffer_bank10_data_29_29_3_lpi_1, buffer_bank10_data_30_29_3_lpi_1,
          buffer_bank10_data_31_29_3_lpi_1, buffer_bank10_data_32_29_3_lpi_1, buffer_bank10_data_33_29_3_lpi_1,
          buffer_bank10_data_34_29_3_lpi_1, buffer_bank10_data_35_29_3_lpi_1, buffer_bank10_data_36_29_3_lpi_1,
          buffer_bank10_data_37_29_3_lpi_1, buffer_bank10_data_38_29_3_lpi_1, buffer_bank10_data_39_29_3_lpi_1,
          buffer_bank10_data_40_29_3_lpi_1, buffer_bank10_data_41_29_3_lpi_1, buffer_bank10_data_42_29_3_lpi_1,
          buffer_bank10_data_43_29_3_lpi_1, buffer_bank10_data_44_29_3_lpi_1, buffer_bank10_data_45_29_3_lpi_1,
          buffer_bank10_data_46_29_3_lpi_1, buffer_bank10_data_47_29_3_lpi_1, buffer_bank10_data_48_29_3_lpi_1,
          buffer_bank10_data_49_29_3_lpi_1, buffer_bank10_data_50_29_3_lpi_1, buffer_bank10_data_51_29_3_lpi_1,
          buffer_bank10_data_52_29_3_lpi_1, buffer_bank10_data_53_29_3_lpi_1, buffer_bank10_data_54_29_3_lpi_1,
          buffer_bank10_data_55_29_3_lpi_1, buffer_bank10_data_56_29_3_lpi_1, buffer_bank10_data_57_29_3_lpi_1,
          buffer_bank10_data_58_29_3_lpi_1, buffer_bank10_data_59_29_3_lpi_1, buffer_bank10_data_60_29_3_lpi_1,
          buffer_bank10_data_61_29_3_lpi_1, buffer_bank10_data_62_29_3_lpi_1, (quads_in_crt_lpi_1[349:323]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_31_24 <= MUX_v_8_64_2(buffer_bank0_data_0_31_24_lpi_1,
          buffer_bank0_data_1_31_24_lpi_1, buffer_bank0_data_2_31_24_lpi_1, buffer_bank0_data_3_31_24_lpi_1,
          buffer_bank0_data_4_31_24_lpi_1, buffer_bank0_data_5_31_24_lpi_1, buffer_bank0_data_6_31_24_lpi_1,
          buffer_bank0_data_7_31_24_lpi_1, buffer_bank0_data_8_31_24_lpi_1, buffer_bank0_data_9_31_24_lpi_1,
          buffer_bank0_data_10_31_24_lpi_1, buffer_bank0_data_11_31_24_lpi_1, buffer_bank0_data_12_31_24_lpi_1,
          buffer_bank0_data_13_31_24_lpi_1, buffer_bank0_data_14_31_24_lpi_1, buffer_bank0_data_15_31_24_lpi_1,
          buffer_bank0_data_16_31_24_lpi_1, buffer_bank0_data_17_31_24_lpi_1, buffer_bank0_data_18_31_24_lpi_1,
          buffer_bank0_data_19_31_24_lpi_1, buffer_bank0_data_20_31_24_lpi_1, buffer_bank0_data_21_31_24_lpi_1,
          buffer_bank0_data_22_31_24_lpi_1, buffer_bank0_data_23_31_24_lpi_1, buffer_bank0_data_24_31_24_lpi_1,
          buffer_bank0_data_25_31_24_lpi_1, buffer_bank0_data_26_31_24_lpi_1, buffer_bank0_data_27_31_24_lpi_1,
          buffer_bank0_data_28_31_24_lpi_1, buffer_bank0_data_29_31_24_lpi_1, buffer_bank0_data_30_31_24_lpi_1,
          buffer_bank0_data_31_31_24_lpi_1, buffer_bank0_data_32_31_24_lpi_1, buffer_bank0_data_33_31_24_lpi_1,
          buffer_bank0_data_34_31_24_lpi_1, buffer_bank0_data_35_31_24_lpi_1, buffer_bank0_data_36_31_24_lpi_1,
          buffer_bank0_data_37_31_24_lpi_1, buffer_bank0_data_38_31_24_lpi_1, buffer_bank0_data_39_31_24_lpi_1,
          buffer_bank0_data_40_31_24_lpi_1, buffer_bank0_data_41_31_24_lpi_1, buffer_bank0_data_42_31_24_lpi_1,
          buffer_bank0_data_43_31_24_lpi_1, buffer_bank0_data_44_31_24_lpi_1, buffer_bank0_data_45_31_24_lpi_1,
          buffer_bank0_data_46_31_24_lpi_1, buffer_bank0_data_47_31_24_lpi_1, buffer_bank0_data_48_31_24_lpi_1,
          buffer_bank0_data_49_31_24_lpi_1, buffer_bank0_data_50_31_24_lpi_1, buffer_bank0_data_51_31_24_lpi_1,
          buffer_bank0_data_52_31_24_lpi_1, buffer_bank0_data_53_31_24_lpi_1, buffer_bank0_data_54_31_24_lpi_1,
          buffer_bank0_data_55_31_24_lpi_1, buffer_bank0_data_56_31_24_lpi_1, buffer_bank0_data_57_31_24_lpi_1,
          buffer_bank0_data_58_31_24_lpi_1, buffer_bank0_data_59_31_24_lpi_1, buffer_bank0_data_60_31_24_lpi_1,
          buffer_bank0_data_61_31_24_lpi_1, buffer_bank0_data_62_31_24_lpi_1, (quads_in_crt_lpi_1[31:24]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_322_320 <= MUX_v_3_64_2(buffer_bank10_data_0_2_0_lpi_1,
          buffer_bank10_data_1_2_0_lpi_1, buffer_bank10_data_2_2_0_lpi_1, buffer_bank10_data_3_2_0_lpi_1,
          buffer_bank10_data_4_2_0_lpi_1, buffer_bank10_data_5_2_0_lpi_1, buffer_bank10_data_6_2_0_lpi_1,
          buffer_bank10_data_7_2_0_lpi_1, buffer_bank10_data_8_2_0_lpi_1, buffer_bank10_data_9_2_0_lpi_1,
          buffer_bank10_data_10_2_0_lpi_1, buffer_bank10_data_11_2_0_lpi_1, buffer_bank10_data_12_2_0_lpi_1,
          buffer_bank10_data_13_2_0_lpi_1, buffer_bank10_data_14_2_0_lpi_1, buffer_bank10_data_15_2_0_lpi_1,
          buffer_bank10_data_16_2_0_lpi_1, buffer_bank10_data_17_2_0_lpi_1, buffer_bank10_data_18_2_0_lpi_1,
          buffer_bank10_data_19_2_0_lpi_1, buffer_bank10_data_20_2_0_lpi_1, buffer_bank10_data_21_2_0_lpi_1,
          buffer_bank10_data_22_2_0_lpi_1, buffer_bank10_data_23_2_0_lpi_1, buffer_bank10_data_24_2_0_lpi_1,
          buffer_bank10_data_25_2_0_lpi_1, buffer_bank10_data_26_2_0_lpi_1, buffer_bank10_data_27_2_0_lpi_1,
          buffer_bank10_data_28_2_0_lpi_1, buffer_bank10_data_29_2_0_lpi_1, buffer_bank10_data_30_2_0_lpi_1,
          buffer_bank10_data_31_2_0_lpi_1, buffer_bank10_data_32_2_0_lpi_1, buffer_bank10_data_33_2_0_lpi_1,
          buffer_bank10_data_34_2_0_lpi_1, buffer_bank10_data_35_2_0_lpi_1, buffer_bank10_data_36_2_0_lpi_1,
          buffer_bank10_data_37_2_0_lpi_1, buffer_bank10_data_38_2_0_lpi_1, buffer_bank10_data_39_2_0_lpi_1,
          buffer_bank10_data_40_2_0_lpi_1, buffer_bank10_data_41_2_0_lpi_1, buffer_bank10_data_42_2_0_lpi_1,
          buffer_bank10_data_43_2_0_lpi_1, buffer_bank10_data_44_2_0_lpi_1, buffer_bank10_data_45_2_0_lpi_1,
          buffer_bank10_data_46_2_0_lpi_1, buffer_bank10_data_47_2_0_lpi_1, buffer_bank10_data_48_2_0_lpi_1,
          buffer_bank10_data_49_2_0_lpi_1, buffer_bank10_data_50_2_0_lpi_1, buffer_bank10_data_51_2_0_lpi_1,
          buffer_bank10_data_52_2_0_lpi_1, buffer_bank10_data_53_2_0_lpi_1, buffer_bank10_data_54_2_0_lpi_1,
          buffer_bank10_data_55_2_0_lpi_1, buffer_bank10_data_56_2_0_lpi_1, buffer_bank10_data_57_2_0_lpi_1,
          buffer_bank10_data_58_2_0_lpi_1, buffer_bank10_data_59_2_0_lpi_1, buffer_bank10_data_60_2_0_lpi_1,
          buffer_bank10_data_61_2_0_lpi_1, buffer_bank10_data_62_2_0_lpi_1, (quads_in_crt_lpi_1[322:320]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_35_32 <= MUX_v_4_64_2(buffer_bank1_data_0_3_0_lpi_1, buffer_bank1_data_1_3_0_lpi_1,
          buffer_bank1_data_2_3_0_lpi_1, buffer_bank1_data_3_3_0_lpi_1, buffer_bank1_data_4_3_0_lpi_1,
          buffer_bank1_data_5_3_0_lpi_1, buffer_bank1_data_6_3_0_lpi_1, buffer_bank1_data_7_3_0_lpi_1,
          buffer_bank1_data_8_3_0_lpi_1, buffer_bank1_data_9_3_0_lpi_1, buffer_bank1_data_10_3_0_lpi_1,
          buffer_bank1_data_11_3_0_lpi_1, buffer_bank1_data_12_3_0_lpi_1, buffer_bank1_data_13_3_0_lpi_1,
          buffer_bank1_data_14_3_0_lpi_1, buffer_bank1_data_15_3_0_lpi_1, buffer_bank1_data_16_3_0_lpi_1,
          buffer_bank1_data_17_3_0_lpi_1, buffer_bank1_data_18_3_0_lpi_1, buffer_bank1_data_19_3_0_lpi_1,
          buffer_bank1_data_20_3_0_lpi_1, buffer_bank1_data_21_3_0_lpi_1, buffer_bank1_data_22_3_0_lpi_1,
          buffer_bank1_data_23_3_0_lpi_1, buffer_bank1_data_24_3_0_lpi_1, buffer_bank1_data_25_3_0_lpi_1,
          buffer_bank1_data_26_3_0_lpi_1, buffer_bank1_data_27_3_0_lpi_1, buffer_bank1_data_28_3_0_lpi_1,
          buffer_bank1_data_29_3_0_lpi_1, buffer_bank1_data_30_3_0_lpi_1, buffer_bank1_data_31_3_0_lpi_1,
          buffer_bank1_data_32_3_0_lpi_1, buffer_bank1_data_33_3_0_lpi_1, buffer_bank1_data_34_3_0_lpi_1,
          buffer_bank1_data_35_3_0_lpi_1, buffer_bank1_data_36_3_0_lpi_1, buffer_bank1_data_37_3_0_lpi_1,
          buffer_bank1_data_38_3_0_lpi_1, buffer_bank1_data_39_3_0_lpi_1, buffer_bank1_data_40_3_0_lpi_1,
          buffer_bank1_data_41_3_0_lpi_1, buffer_bank1_data_42_3_0_lpi_1, buffer_bank1_data_43_3_0_lpi_1,
          buffer_bank1_data_44_3_0_lpi_1, buffer_bank1_data_45_3_0_lpi_1, buffer_bank1_data_46_3_0_lpi_1,
          buffer_bank1_data_47_3_0_lpi_1, buffer_bank1_data_48_3_0_lpi_1, buffer_bank1_data_49_3_0_lpi_1,
          buffer_bank1_data_50_3_0_lpi_1, buffer_bank1_data_51_3_0_lpi_1, buffer_bank1_data_52_3_0_lpi_1,
          buffer_bank1_data_53_3_0_lpi_1, buffer_bank1_data_54_3_0_lpi_1, buffer_bank1_data_55_3_0_lpi_1,
          buffer_bank1_data_56_3_0_lpi_1, buffer_bank1_data_57_3_0_lpi_1, buffer_bank1_data_58_3_0_lpi_1,
          buffer_bank1_data_59_3_0_lpi_1, buffer_bank1_data_60_3_0_lpi_1, buffer_bank1_data_61_3_0_lpi_1,
          buffer_bank1_data_62_3_0_lpi_1, (quads_in_crt_lpi_1[35:32]), for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_319_296 <= MUX_v_24_64_2(buffer_bank9_data_0_31_8_lpi_1,
          buffer_bank9_data_1_31_8_lpi_1, buffer_bank9_data_2_31_8_lpi_1, buffer_bank9_data_3_31_8_lpi_1,
          buffer_bank9_data_4_31_8_lpi_1, buffer_bank9_data_5_31_8_lpi_1, buffer_bank9_data_6_31_8_lpi_1,
          buffer_bank9_data_7_31_8_lpi_1, buffer_bank9_data_8_31_8_lpi_1, buffer_bank9_data_9_31_8_lpi_1,
          buffer_bank9_data_10_31_8_lpi_1, buffer_bank9_data_11_31_8_lpi_1, buffer_bank9_data_12_31_8_lpi_1,
          buffer_bank9_data_13_31_8_lpi_1, buffer_bank9_data_14_31_8_lpi_1, buffer_bank9_data_15_31_8_lpi_1,
          buffer_bank9_data_16_31_8_lpi_1, buffer_bank9_data_17_31_8_lpi_1, buffer_bank9_data_18_31_8_lpi_1,
          buffer_bank9_data_19_31_8_lpi_1, buffer_bank9_data_20_31_8_lpi_1, buffer_bank9_data_21_31_8_lpi_1,
          buffer_bank9_data_22_31_8_lpi_1, buffer_bank9_data_23_31_8_lpi_1, buffer_bank9_data_24_31_8_lpi_1,
          buffer_bank9_data_25_31_8_lpi_1, buffer_bank9_data_26_31_8_lpi_1, buffer_bank9_data_27_31_8_lpi_1,
          buffer_bank9_data_28_31_8_lpi_1, buffer_bank9_data_29_31_8_lpi_1, buffer_bank9_data_30_31_8_lpi_1,
          buffer_bank9_data_31_31_8_lpi_1, buffer_bank9_data_32_31_8_lpi_1, buffer_bank9_data_33_31_8_lpi_1,
          buffer_bank9_data_34_31_8_lpi_1, buffer_bank9_data_35_31_8_lpi_1, buffer_bank9_data_36_31_8_lpi_1,
          buffer_bank9_data_37_31_8_lpi_1, buffer_bank9_data_38_31_8_lpi_1, buffer_bank9_data_39_31_8_lpi_1,
          buffer_bank9_data_40_31_8_lpi_1, buffer_bank9_data_41_31_8_lpi_1, buffer_bank9_data_42_31_8_lpi_1,
          buffer_bank9_data_43_31_8_lpi_1, buffer_bank9_data_44_31_8_lpi_1, buffer_bank9_data_45_31_8_lpi_1,
          buffer_bank9_data_46_31_8_lpi_1, buffer_bank9_data_47_31_8_lpi_1, buffer_bank9_data_48_31_8_lpi_1,
          buffer_bank9_data_49_31_8_lpi_1, buffer_bank9_data_50_31_8_lpi_1, buffer_bank9_data_51_31_8_lpi_1,
          buffer_bank9_data_52_31_8_lpi_1, buffer_bank9_data_53_31_8_lpi_1, buffer_bank9_data_54_31_8_lpi_1,
          buffer_bank9_data_55_31_8_lpi_1, buffer_bank9_data_56_31_8_lpi_1, buffer_bank9_data_57_31_8_lpi_1,
          buffer_bank9_data_58_31_8_lpi_1, buffer_bank9_data_59_31_8_lpi_1, buffer_bank9_data_60_31_8_lpi_1,
          buffer_bank9_data_61_31_8_lpi_1, buffer_bank9_data_62_31_8_lpi_1, (quads_in_crt_lpi_1[319:296]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_47_36 <= MUX_v_12_64_2(buffer_bank1_data_0_15_4_lpi_1,
          buffer_bank1_data_1_15_4_lpi_1, buffer_bank1_data_2_15_4_lpi_1, buffer_bank1_data_3_15_4_lpi_1,
          buffer_bank1_data_4_15_4_lpi_1, buffer_bank1_data_5_15_4_lpi_1, buffer_bank1_data_6_15_4_lpi_1,
          buffer_bank1_data_7_15_4_lpi_1, buffer_bank1_data_8_15_4_lpi_1, buffer_bank1_data_9_15_4_lpi_1,
          buffer_bank1_data_10_15_4_lpi_1, buffer_bank1_data_11_15_4_lpi_1, buffer_bank1_data_12_15_4_lpi_1,
          buffer_bank1_data_13_15_4_lpi_1, buffer_bank1_data_14_15_4_lpi_1, buffer_bank1_data_15_15_4_lpi_1,
          buffer_bank1_data_16_15_4_lpi_1, buffer_bank1_data_17_15_4_lpi_1, buffer_bank1_data_18_15_4_lpi_1,
          buffer_bank1_data_19_15_4_lpi_1, buffer_bank1_data_20_15_4_lpi_1, buffer_bank1_data_21_15_4_lpi_1,
          buffer_bank1_data_22_15_4_lpi_1, buffer_bank1_data_23_15_4_lpi_1, buffer_bank1_data_24_15_4_lpi_1,
          buffer_bank1_data_25_15_4_lpi_1, buffer_bank1_data_26_15_4_lpi_1, buffer_bank1_data_27_15_4_lpi_1,
          buffer_bank1_data_28_15_4_lpi_1, buffer_bank1_data_29_15_4_lpi_1, buffer_bank1_data_30_15_4_lpi_1,
          buffer_bank1_data_31_15_4_lpi_1, buffer_bank1_data_32_15_4_lpi_1, buffer_bank1_data_33_15_4_lpi_1,
          buffer_bank1_data_34_15_4_lpi_1, buffer_bank1_data_35_15_4_lpi_1, buffer_bank1_data_36_15_4_lpi_1,
          buffer_bank1_data_37_15_4_lpi_1, buffer_bank1_data_38_15_4_lpi_1, buffer_bank1_data_39_15_4_lpi_1,
          buffer_bank1_data_40_15_4_lpi_1, buffer_bank1_data_41_15_4_lpi_1, buffer_bank1_data_42_15_4_lpi_1,
          buffer_bank1_data_43_15_4_lpi_1, buffer_bank1_data_44_15_4_lpi_1, buffer_bank1_data_45_15_4_lpi_1,
          buffer_bank1_data_46_15_4_lpi_1, buffer_bank1_data_47_15_4_lpi_1, buffer_bank1_data_48_15_4_lpi_1,
          buffer_bank1_data_49_15_4_lpi_1, buffer_bank1_data_50_15_4_lpi_1, buffer_bank1_data_51_15_4_lpi_1,
          buffer_bank1_data_52_15_4_lpi_1, buffer_bank1_data_53_15_4_lpi_1, buffer_bank1_data_54_15_4_lpi_1,
          buffer_bank1_data_55_15_4_lpi_1, buffer_bank1_data_56_15_4_lpi_1, buffer_bank1_data_57_15_4_lpi_1,
          buffer_bank1_data_58_15_4_lpi_1, buffer_bank1_data_59_15_4_lpi_1, buffer_bank1_data_60_15_4_lpi_1,
          buffer_bank1_data_61_15_4_lpi_1, buffer_bank1_data_62_15_4_lpi_1, (quads_in_crt_lpi_1[47:36]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_295_288 <= MUX_v_8_64_2(buffer_bank9_data_0_7_0_lpi_1,
          buffer_bank9_data_1_7_0_lpi_1, buffer_bank9_data_2_7_0_lpi_1, buffer_bank9_data_3_7_0_lpi_1,
          buffer_bank9_data_4_7_0_lpi_1, buffer_bank9_data_5_7_0_lpi_1, buffer_bank9_data_6_7_0_lpi_1,
          buffer_bank9_data_7_7_0_lpi_1, buffer_bank9_data_8_7_0_lpi_1, buffer_bank9_data_9_7_0_lpi_1,
          buffer_bank9_data_10_7_0_lpi_1, buffer_bank9_data_11_7_0_lpi_1, buffer_bank9_data_12_7_0_lpi_1,
          buffer_bank9_data_13_7_0_lpi_1, buffer_bank9_data_14_7_0_lpi_1, buffer_bank9_data_15_7_0_lpi_1,
          buffer_bank9_data_16_7_0_lpi_1, buffer_bank9_data_17_7_0_lpi_1, buffer_bank9_data_18_7_0_lpi_1,
          buffer_bank9_data_19_7_0_lpi_1, buffer_bank9_data_20_7_0_lpi_1, buffer_bank9_data_21_7_0_lpi_1,
          buffer_bank9_data_22_7_0_lpi_1, buffer_bank9_data_23_7_0_lpi_1, buffer_bank9_data_24_7_0_lpi_1,
          buffer_bank9_data_25_7_0_lpi_1, buffer_bank9_data_26_7_0_lpi_1, buffer_bank9_data_27_7_0_lpi_1,
          buffer_bank9_data_28_7_0_lpi_1, buffer_bank9_data_29_7_0_lpi_1, buffer_bank9_data_30_7_0_lpi_1,
          buffer_bank9_data_31_7_0_lpi_1, buffer_bank9_data_32_7_0_lpi_1, buffer_bank9_data_33_7_0_lpi_1,
          buffer_bank9_data_34_7_0_lpi_1, buffer_bank9_data_35_7_0_lpi_1, buffer_bank9_data_36_7_0_lpi_1,
          buffer_bank9_data_37_7_0_lpi_1, buffer_bank9_data_38_7_0_lpi_1, buffer_bank9_data_39_7_0_lpi_1,
          buffer_bank9_data_40_7_0_lpi_1, buffer_bank9_data_41_7_0_lpi_1, buffer_bank9_data_42_7_0_lpi_1,
          buffer_bank9_data_43_7_0_lpi_1, buffer_bank9_data_44_7_0_lpi_1, buffer_bank9_data_45_7_0_lpi_1,
          buffer_bank9_data_46_7_0_lpi_1, buffer_bank9_data_47_7_0_lpi_1, buffer_bank9_data_48_7_0_lpi_1,
          buffer_bank9_data_49_7_0_lpi_1, buffer_bank9_data_50_7_0_lpi_1, buffer_bank9_data_51_7_0_lpi_1,
          buffer_bank9_data_52_7_0_lpi_1, buffer_bank9_data_53_7_0_lpi_1, buffer_bank9_data_54_7_0_lpi_1,
          buffer_bank9_data_55_7_0_lpi_1, buffer_bank9_data_56_7_0_lpi_1, buffer_bank9_data_57_7_0_lpi_1,
          buffer_bank9_data_58_7_0_lpi_1, buffer_bank9_data_59_7_0_lpi_1, buffer_bank9_data_60_7_0_lpi_1,
          buffer_bank9_data_61_7_0_lpi_1, buffer_bank9_data_62_7_0_lpi_1, (quads_in_crt_lpi_1[295:288]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_59_48 <= MUX_v_12_64_2(buffer_bank1_data_0_27_16_lpi_1,
          buffer_bank1_data_1_27_16_lpi_1, buffer_bank1_data_2_27_16_lpi_1, buffer_bank1_data_3_27_16_lpi_1,
          buffer_bank1_data_4_27_16_lpi_1, buffer_bank1_data_5_27_16_lpi_1, buffer_bank1_data_6_27_16_lpi_1,
          buffer_bank1_data_7_27_16_lpi_1, buffer_bank1_data_8_27_16_lpi_1, buffer_bank1_data_9_27_16_lpi_1,
          buffer_bank1_data_10_27_16_lpi_1, buffer_bank1_data_11_27_16_lpi_1, buffer_bank1_data_12_27_16_lpi_1,
          buffer_bank1_data_13_27_16_lpi_1, buffer_bank1_data_14_27_16_lpi_1, buffer_bank1_data_15_27_16_lpi_1,
          buffer_bank1_data_16_27_16_lpi_1, buffer_bank1_data_17_27_16_lpi_1, buffer_bank1_data_18_27_16_lpi_1,
          buffer_bank1_data_19_27_16_lpi_1, buffer_bank1_data_20_27_16_lpi_1, buffer_bank1_data_21_27_16_lpi_1,
          buffer_bank1_data_22_27_16_lpi_1, buffer_bank1_data_23_27_16_lpi_1, buffer_bank1_data_24_27_16_lpi_1,
          buffer_bank1_data_25_27_16_lpi_1, buffer_bank1_data_26_27_16_lpi_1, buffer_bank1_data_27_27_16_lpi_1,
          buffer_bank1_data_28_27_16_lpi_1, buffer_bank1_data_29_27_16_lpi_1, buffer_bank1_data_30_27_16_lpi_1,
          buffer_bank1_data_31_27_16_lpi_1, buffer_bank1_data_32_27_16_lpi_1, buffer_bank1_data_33_27_16_lpi_1,
          buffer_bank1_data_34_27_16_lpi_1, buffer_bank1_data_35_27_16_lpi_1, buffer_bank1_data_36_27_16_lpi_1,
          buffer_bank1_data_37_27_16_lpi_1, buffer_bank1_data_38_27_16_lpi_1, buffer_bank1_data_39_27_16_lpi_1,
          buffer_bank1_data_40_27_16_lpi_1, buffer_bank1_data_41_27_16_lpi_1, buffer_bank1_data_42_27_16_lpi_1,
          buffer_bank1_data_43_27_16_lpi_1, buffer_bank1_data_44_27_16_lpi_1, buffer_bank1_data_45_27_16_lpi_1,
          buffer_bank1_data_46_27_16_lpi_1, buffer_bank1_data_47_27_16_lpi_1, buffer_bank1_data_48_27_16_lpi_1,
          buffer_bank1_data_49_27_16_lpi_1, buffer_bank1_data_50_27_16_lpi_1, buffer_bank1_data_51_27_16_lpi_1,
          buffer_bank1_data_52_27_16_lpi_1, buffer_bank1_data_53_27_16_lpi_1, buffer_bank1_data_54_27_16_lpi_1,
          buffer_bank1_data_55_27_16_lpi_1, buffer_bank1_data_56_27_16_lpi_1, buffer_bank1_data_57_27_16_lpi_1,
          buffer_bank1_data_58_27_16_lpi_1, buffer_bank1_data_59_27_16_lpi_1, buffer_bank1_data_60_27_16_lpi_1,
          buffer_bank1_data_61_27_16_lpi_1, buffer_bank1_data_62_27_16_lpi_1, (quads_in_crt_lpi_1[59:48]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_287_265 <= MUX_v_23_64_2(buffer_bank8_data_0_31_9_lpi_1,
          buffer_bank8_data_1_31_9_lpi_1, buffer_bank8_data_2_31_9_lpi_1, buffer_bank8_data_3_31_9_lpi_1,
          buffer_bank8_data_4_31_9_lpi_1, buffer_bank8_data_5_31_9_lpi_1, buffer_bank8_data_6_31_9_lpi_1,
          buffer_bank8_data_7_31_9_lpi_1, buffer_bank8_data_8_31_9_lpi_1, buffer_bank8_data_9_31_9_lpi_1,
          buffer_bank8_data_10_31_9_lpi_1, buffer_bank8_data_11_31_9_lpi_1, buffer_bank8_data_12_31_9_lpi_1,
          buffer_bank8_data_13_31_9_lpi_1, buffer_bank8_data_14_31_9_lpi_1, buffer_bank8_data_15_31_9_lpi_1,
          buffer_bank8_data_16_31_9_lpi_1, buffer_bank8_data_17_31_9_lpi_1, buffer_bank8_data_18_31_9_lpi_1,
          buffer_bank8_data_19_31_9_lpi_1, buffer_bank8_data_20_31_9_lpi_1, buffer_bank8_data_21_31_9_lpi_1,
          buffer_bank8_data_22_31_9_lpi_1, buffer_bank8_data_23_31_9_lpi_1, buffer_bank8_data_24_31_9_lpi_1,
          buffer_bank8_data_25_31_9_lpi_1, buffer_bank8_data_26_31_9_lpi_1, buffer_bank8_data_27_31_9_lpi_1,
          buffer_bank8_data_28_31_9_lpi_1, buffer_bank8_data_29_31_9_lpi_1, buffer_bank8_data_30_31_9_lpi_1,
          buffer_bank8_data_31_31_9_lpi_1, buffer_bank8_data_32_31_9_lpi_1, buffer_bank8_data_33_31_9_lpi_1,
          buffer_bank8_data_34_31_9_lpi_1, buffer_bank8_data_35_31_9_lpi_1, buffer_bank8_data_36_31_9_lpi_1,
          buffer_bank8_data_37_31_9_lpi_1, buffer_bank8_data_38_31_9_lpi_1, buffer_bank8_data_39_31_9_lpi_1,
          buffer_bank8_data_40_31_9_lpi_1, buffer_bank8_data_41_31_9_lpi_1, buffer_bank8_data_42_31_9_lpi_1,
          buffer_bank8_data_43_31_9_lpi_1, buffer_bank8_data_44_31_9_lpi_1, buffer_bank8_data_45_31_9_lpi_1,
          buffer_bank8_data_46_31_9_lpi_1, buffer_bank8_data_47_31_9_lpi_1, buffer_bank8_data_48_31_9_lpi_1,
          buffer_bank8_data_49_31_9_lpi_1, buffer_bank8_data_50_31_9_lpi_1, buffer_bank8_data_51_31_9_lpi_1,
          buffer_bank8_data_52_31_9_lpi_1, buffer_bank8_data_53_31_9_lpi_1, buffer_bank8_data_54_31_9_lpi_1,
          buffer_bank8_data_55_31_9_lpi_1, buffer_bank8_data_56_31_9_lpi_1, buffer_bank8_data_57_31_9_lpi_1,
          buffer_bank8_data_58_31_9_lpi_1, buffer_bank8_data_59_31_9_lpi_1, buffer_bank8_data_60_31_9_lpi_1,
          buffer_bank8_data_61_31_9_lpi_1, buffer_bank8_data_62_31_9_lpi_1, (quads_in_crt_lpi_1[287:265]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_63_60 <= MUX_v_4_64_2(buffer_bank1_data_0_31_28_lpi_1,
          buffer_bank1_data_1_31_28_lpi_1, buffer_bank1_data_2_31_28_lpi_1, buffer_bank1_data_3_31_28_lpi_1,
          buffer_bank1_data_4_31_28_lpi_1, buffer_bank1_data_5_31_28_lpi_1, buffer_bank1_data_6_31_28_lpi_1,
          buffer_bank1_data_7_31_28_lpi_1, buffer_bank1_data_8_31_28_lpi_1, buffer_bank1_data_9_31_28_lpi_1,
          buffer_bank1_data_10_31_28_lpi_1, buffer_bank1_data_11_31_28_lpi_1, buffer_bank1_data_12_31_28_lpi_1,
          buffer_bank1_data_13_31_28_lpi_1, buffer_bank1_data_14_31_28_lpi_1, buffer_bank1_data_15_31_28_lpi_1,
          buffer_bank1_data_16_31_28_lpi_1, buffer_bank1_data_17_31_28_lpi_1, buffer_bank1_data_18_31_28_lpi_1,
          buffer_bank1_data_19_31_28_lpi_1, buffer_bank1_data_20_31_28_lpi_1, buffer_bank1_data_21_31_28_lpi_1,
          buffer_bank1_data_22_31_28_lpi_1, buffer_bank1_data_23_31_28_lpi_1, buffer_bank1_data_24_31_28_lpi_1,
          buffer_bank1_data_25_31_28_lpi_1, buffer_bank1_data_26_31_28_lpi_1, buffer_bank1_data_27_31_28_lpi_1,
          buffer_bank1_data_28_31_28_lpi_1, buffer_bank1_data_29_31_28_lpi_1, buffer_bank1_data_30_31_28_lpi_1,
          buffer_bank1_data_31_31_28_lpi_1, buffer_bank1_data_32_31_28_lpi_1, buffer_bank1_data_33_31_28_lpi_1,
          buffer_bank1_data_34_31_28_lpi_1, buffer_bank1_data_35_31_28_lpi_1, buffer_bank1_data_36_31_28_lpi_1,
          buffer_bank1_data_37_31_28_lpi_1, buffer_bank1_data_38_31_28_lpi_1, buffer_bank1_data_39_31_28_lpi_1,
          buffer_bank1_data_40_31_28_lpi_1, buffer_bank1_data_41_31_28_lpi_1, buffer_bank1_data_42_31_28_lpi_1,
          buffer_bank1_data_43_31_28_lpi_1, buffer_bank1_data_44_31_28_lpi_1, buffer_bank1_data_45_31_28_lpi_1,
          buffer_bank1_data_46_31_28_lpi_1, buffer_bank1_data_47_31_28_lpi_1, buffer_bank1_data_48_31_28_lpi_1,
          buffer_bank1_data_49_31_28_lpi_1, buffer_bank1_data_50_31_28_lpi_1, buffer_bank1_data_51_31_28_lpi_1,
          buffer_bank1_data_52_31_28_lpi_1, buffer_bank1_data_53_31_28_lpi_1, buffer_bank1_data_54_31_28_lpi_1,
          buffer_bank1_data_55_31_28_lpi_1, buffer_bank1_data_56_31_28_lpi_1, buffer_bank1_data_57_31_28_lpi_1,
          buffer_bank1_data_58_31_28_lpi_1, buffer_bank1_data_59_31_28_lpi_1, buffer_bank1_data_60_31_28_lpi_1,
          buffer_bank1_data_61_31_28_lpi_1, buffer_bank1_data_62_31_28_lpi_1, (quads_in_crt_lpi_1[63:60]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_264_256 <= MUX_v_9_64_2(buffer_bank8_data_0_8_0_lpi_1,
          buffer_bank8_data_1_8_0_lpi_1, buffer_bank8_data_2_8_0_lpi_1, buffer_bank8_data_3_8_0_lpi_1,
          buffer_bank8_data_4_8_0_lpi_1, buffer_bank8_data_5_8_0_lpi_1, buffer_bank8_data_6_8_0_lpi_1,
          buffer_bank8_data_7_8_0_lpi_1, buffer_bank8_data_8_8_0_lpi_1, buffer_bank8_data_9_8_0_lpi_1,
          buffer_bank8_data_10_8_0_lpi_1, buffer_bank8_data_11_8_0_lpi_1, buffer_bank8_data_12_8_0_lpi_1,
          buffer_bank8_data_13_8_0_lpi_1, buffer_bank8_data_14_8_0_lpi_1, buffer_bank8_data_15_8_0_lpi_1,
          buffer_bank8_data_16_8_0_lpi_1, buffer_bank8_data_17_8_0_lpi_1, buffer_bank8_data_18_8_0_lpi_1,
          buffer_bank8_data_19_8_0_lpi_1, buffer_bank8_data_20_8_0_lpi_1, buffer_bank8_data_21_8_0_lpi_1,
          buffer_bank8_data_22_8_0_lpi_1, buffer_bank8_data_23_8_0_lpi_1, buffer_bank8_data_24_8_0_lpi_1,
          buffer_bank8_data_25_8_0_lpi_1, buffer_bank8_data_26_8_0_lpi_1, buffer_bank8_data_27_8_0_lpi_1,
          buffer_bank8_data_28_8_0_lpi_1, buffer_bank8_data_29_8_0_lpi_1, buffer_bank8_data_30_8_0_lpi_1,
          buffer_bank8_data_31_8_0_lpi_1, buffer_bank8_data_32_8_0_lpi_1, buffer_bank8_data_33_8_0_lpi_1,
          buffer_bank8_data_34_8_0_lpi_1, buffer_bank8_data_35_8_0_lpi_1, buffer_bank8_data_36_8_0_lpi_1,
          buffer_bank8_data_37_8_0_lpi_1, buffer_bank8_data_38_8_0_lpi_1, buffer_bank8_data_39_8_0_lpi_1,
          buffer_bank8_data_40_8_0_lpi_1, buffer_bank8_data_41_8_0_lpi_1, buffer_bank8_data_42_8_0_lpi_1,
          buffer_bank8_data_43_8_0_lpi_1, buffer_bank8_data_44_8_0_lpi_1, buffer_bank8_data_45_8_0_lpi_1,
          buffer_bank8_data_46_8_0_lpi_1, buffer_bank8_data_47_8_0_lpi_1, buffer_bank8_data_48_8_0_lpi_1,
          buffer_bank8_data_49_8_0_lpi_1, buffer_bank8_data_50_8_0_lpi_1, buffer_bank8_data_51_8_0_lpi_1,
          buffer_bank8_data_52_8_0_lpi_1, buffer_bank8_data_53_8_0_lpi_1, buffer_bank8_data_54_8_0_lpi_1,
          buffer_bank8_data_55_8_0_lpi_1, buffer_bank8_data_56_8_0_lpi_1, buffer_bank8_data_57_8_0_lpi_1,
          buffer_bank8_data_58_8_0_lpi_1, buffer_bank8_data_59_8_0_lpi_1, buffer_bank8_data_60_8_0_lpi_1,
          buffer_bank8_data_61_8_0_lpi_1, buffer_bank8_data_62_8_0_lpi_1, (quads_in_crt_lpi_1[264:256]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_71_64 <= MUX_v_8_64_2(buffer_bank2_data_0_7_0_lpi_1, buffer_bank2_data_1_7_0_lpi_1,
          buffer_bank2_data_2_7_0_lpi_1, buffer_bank2_data_3_7_0_lpi_1, buffer_bank2_data_4_7_0_lpi_1,
          buffer_bank2_data_5_7_0_lpi_1, buffer_bank2_data_6_7_0_lpi_1, buffer_bank2_data_7_7_0_lpi_1,
          buffer_bank2_data_8_7_0_lpi_1, buffer_bank2_data_9_7_0_lpi_1, buffer_bank2_data_10_7_0_lpi_1,
          buffer_bank2_data_11_7_0_lpi_1, buffer_bank2_data_12_7_0_lpi_1, buffer_bank2_data_13_7_0_lpi_1,
          buffer_bank2_data_14_7_0_lpi_1, buffer_bank2_data_15_7_0_lpi_1, buffer_bank2_data_16_7_0_lpi_1,
          buffer_bank2_data_17_7_0_lpi_1, buffer_bank2_data_18_7_0_lpi_1, buffer_bank2_data_19_7_0_lpi_1,
          buffer_bank2_data_20_7_0_lpi_1, buffer_bank2_data_21_7_0_lpi_1, buffer_bank2_data_22_7_0_lpi_1,
          buffer_bank2_data_23_7_0_lpi_1, buffer_bank2_data_24_7_0_lpi_1, buffer_bank2_data_25_7_0_lpi_1,
          buffer_bank2_data_26_7_0_lpi_1, buffer_bank2_data_27_7_0_lpi_1, buffer_bank2_data_28_7_0_lpi_1,
          buffer_bank2_data_29_7_0_lpi_1, buffer_bank2_data_30_7_0_lpi_1, buffer_bank2_data_31_7_0_lpi_1,
          buffer_bank2_data_32_7_0_lpi_1, buffer_bank2_data_33_7_0_lpi_1, buffer_bank2_data_34_7_0_lpi_1,
          buffer_bank2_data_35_7_0_lpi_1, buffer_bank2_data_36_7_0_lpi_1, buffer_bank2_data_37_7_0_lpi_1,
          buffer_bank2_data_38_7_0_lpi_1, buffer_bank2_data_39_7_0_lpi_1, buffer_bank2_data_40_7_0_lpi_1,
          buffer_bank2_data_41_7_0_lpi_1, buffer_bank2_data_42_7_0_lpi_1, buffer_bank2_data_43_7_0_lpi_1,
          buffer_bank2_data_44_7_0_lpi_1, buffer_bank2_data_45_7_0_lpi_1, buffer_bank2_data_46_7_0_lpi_1,
          buffer_bank2_data_47_7_0_lpi_1, buffer_bank2_data_48_7_0_lpi_1, buffer_bank2_data_49_7_0_lpi_1,
          buffer_bank2_data_50_7_0_lpi_1, buffer_bank2_data_51_7_0_lpi_1, buffer_bank2_data_52_7_0_lpi_1,
          buffer_bank2_data_53_7_0_lpi_1, buffer_bank2_data_54_7_0_lpi_1, buffer_bank2_data_55_7_0_lpi_1,
          buffer_bank2_data_56_7_0_lpi_1, buffer_bank2_data_57_7_0_lpi_1, buffer_bank2_data_58_7_0_lpi_1,
          buffer_bank2_data_59_7_0_lpi_1, buffer_bank2_data_60_7_0_lpi_1, buffer_bank2_data_61_7_0_lpi_1,
          buffer_bank2_data_62_7_0_lpi_1, (quads_in_crt_lpi_1[71:64]), for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_255_240 <= MUX_v_16_64_2(buffer_bank7_data_0_31_16_lpi_1,
          buffer_bank7_data_1_31_16_lpi_1, buffer_bank7_data_2_31_16_lpi_1, buffer_bank7_data_3_31_16_lpi_1,
          buffer_bank7_data_4_31_16_lpi_1, buffer_bank7_data_5_31_16_lpi_1, buffer_bank7_data_6_31_16_lpi_1,
          buffer_bank7_data_7_31_16_lpi_1, buffer_bank7_data_8_31_16_lpi_1, buffer_bank7_data_9_31_16_lpi_1,
          buffer_bank7_data_10_31_16_lpi_1, buffer_bank7_data_11_31_16_lpi_1, buffer_bank7_data_12_31_16_lpi_1,
          buffer_bank7_data_13_31_16_lpi_1, buffer_bank7_data_14_31_16_lpi_1, buffer_bank7_data_15_31_16_lpi_1,
          buffer_bank7_data_16_31_16_lpi_1, buffer_bank7_data_17_31_16_lpi_1, buffer_bank7_data_18_31_16_lpi_1,
          buffer_bank7_data_19_31_16_lpi_1, buffer_bank7_data_20_31_16_lpi_1, buffer_bank7_data_21_31_16_lpi_1,
          buffer_bank7_data_22_31_16_lpi_1, buffer_bank7_data_23_31_16_lpi_1, buffer_bank7_data_24_31_16_lpi_1,
          buffer_bank7_data_25_31_16_lpi_1, buffer_bank7_data_26_31_16_lpi_1, buffer_bank7_data_27_31_16_lpi_1,
          buffer_bank7_data_28_31_16_lpi_1, buffer_bank7_data_29_31_16_lpi_1, buffer_bank7_data_30_31_16_lpi_1,
          buffer_bank7_data_31_31_16_lpi_1, buffer_bank7_data_32_31_16_lpi_1, buffer_bank7_data_33_31_16_lpi_1,
          buffer_bank7_data_34_31_16_lpi_1, buffer_bank7_data_35_31_16_lpi_1, buffer_bank7_data_36_31_16_lpi_1,
          buffer_bank7_data_37_31_16_lpi_1, buffer_bank7_data_38_31_16_lpi_1, buffer_bank7_data_39_31_16_lpi_1,
          buffer_bank7_data_40_31_16_lpi_1, buffer_bank7_data_41_31_16_lpi_1, buffer_bank7_data_42_31_16_lpi_1,
          buffer_bank7_data_43_31_16_lpi_1, buffer_bank7_data_44_31_16_lpi_1, buffer_bank7_data_45_31_16_lpi_1,
          buffer_bank7_data_46_31_16_lpi_1, buffer_bank7_data_47_31_16_lpi_1, buffer_bank7_data_48_31_16_lpi_1,
          buffer_bank7_data_49_31_16_lpi_1, buffer_bank7_data_50_31_16_lpi_1, buffer_bank7_data_51_31_16_lpi_1,
          buffer_bank7_data_52_31_16_lpi_1, buffer_bank7_data_53_31_16_lpi_1, buffer_bank7_data_54_31_16_lpi_1,
          buffer_bank7_data_55_31_16_lpi_1, buffer_bank7_data_56_31_16_lpi_1, buffer_bank7_data_57_31_16_lpi_1,
          buffer_bank7_data_58_31_16_lpi_1, buffer_bank7_data_59_31_16_lpi_1, buffer_bank7_data_60_31_16_lpi_1,
          buffer_bank7_data_61_31_16_lpi_1, buffer_bank7_data_62_31_16_lpi_1, (quads_in_crt_lpi_1[255:240]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_83_72 <= MUX_v_12_64_2(buffer_bank2_data_0_19_8_lpi_1,
          buffer_bank2_data_1_19_8_lpi_1, buffer_bank2_data_2_19_8_lpi_1, buffer_bank2_data_3_19_8_lpi_1,
          buffer_bank2_data_4_19_8_lpi_1, buffer_bank2_data_5_19_8_lpi_1, buffer_bank2_data_6_19_8_lpi_1,
          buffer_bank2_data_7_19_8_lpi_1, buffer_bank2_data_8_19_8_lpi_1, buffer_bank2_data_9_19_8_lpi_1,
          buffer_bank2_data_10_19_8_lpi_1, buffer_bank2_data_11_19_8_lpi_1, buffer_bank2_data_12_19_8_lpi_1,
          buffer_bank2_data_13_19_8_lpi_1, buffer_bank2_data_14_19_8_lpi_1, buffer_bank2_data_15_19_8_lpi_1,
          buffer_bank2_data_16_19_8_lpi_1, buffer_bank2_data_17_19_8_lpi_1, buffer_bank2_data_18_19_8_lpi_1,
          buffer_bank2_data_19_19_8_lpi_1, buffer_bank2_data_20_19_8_lpi_1, buffer_bank2_data_21_19_8_lpi_1,
          buffer_bank2_data_22_19_8_lpi_1, buffer_bank2_data_23_19_8_lpi_1, buffer_bank2_data_24_19_8_lpi_1,
          buffer_bank2_data_25_19_8_lpi_1, buffer_bank2_data_26_19_8_lpi_1, buffer_bank2_data_27_19_8_lpi_1,
          buffer_bank2_data_28_19_8_lpi_1, buffer_bank2_data_29_19_8_lpi_1, buffer_bank2_data_30_19_8_lpi_1,
          buffer_bank2_data_31_19_8_lpi_1, buffer_bank2_data_32_19_8_lpi_1, buffer_bank2_data_33_19_8_lpi_1,
          buffer_bank2_data_34_19_8_lpi_1, buffer_bank2_data_35_19_8_lpi_1, buffer_bank2_data_36_19_8_lpi_1,
          buffer_bank2_data_37_19_8_lpi_1, buffer_bank2_data_38_19_8_lpi_1, buffer_bank2_data_39_19_8_lpi_1,
          buffer_bank2_data_40_19_8_lpi_1, buffer_bank2_data_41_19_8_lpi_1, buffer_bank2_data_42_19_8_lpi_1,
          buffer_bank2_data_43_19_8_lpi_1, buffer_bank2_data_44_19_8_lpi_1, buffer_bank2_data_45_19_8_lpi_1,
          buffer_bank2_data_46_19_8_lpi_1, buffer_bank2_data_47_19_8_lpi_1, buffer_bank2_data_48_19_8_lpi_1,
          buffer_bank2_data_49_19_8_lpi_1, buffer_bank2_data_50_19_8_lpi_1, buffer_bank2_data_51_19_8_lpi_1,
          buffer_bank2_data_52_19_8_lpi_1, buffer_bank2_data_53_19_8_lpi_1, buffer_bank2_data_54_19_8_lpi_1,
          buffer_bank2_data_55_19_8_lpi_1, buffer_bank2_data_56_19_8_lpi_1, buffer_bank2_data_57_19_8_lpi_1,
          buffer_bank2_data_58_19_8_lpi_1, buffer_bank2_data_59_19_8_lpi_1, buffer_bank2_data_60_19_8_lpi_1,
          buffer_bank2_data_61_19_8_lpi_1, buffer_bank2_data_62_19_8_lpi_1, (quads_in_crt_lpi_1[83:72]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_239_224 <= MUX_v_16_64_2(buffer_bank7_data_0_15_0_lpi_1,
          buffer_bank7_data_1_15_0_lpi_1, buffer_bank7_data_2_15_0_lpi_1, buffer_bank7_data_3_15_0_lpi_1,
          buffer_bank7_data_4_15_0_lpi_1, buffer_bank7_data_5_15_0_lpi_1, buffer_bank7_data_6_15_0_lpi_1,
          buffer_bank7_data_7_15_0_lpi_1, buffer_bank7_data_8_15_0_lpi_1, buffer_bank7_data_9_15_0_lpi_1,
          buffer_bank7_data_10_15_0_lpi_1, buffer_bank7_data_11_15_0_lpi_1, buffer_bank7_data_12_15_0_lpi_1,
          buffer_bank7_data_13_15_0_lpi_1, buffer_bank7_data_14_15_0_lpi_1, buffer_bank7_data_15_15_0_lpi_1,
          buffer_bank7_data_16_15_0_lpi_1, buffer_bank7_data_17_15_0_lpi_1, buffer_bank7_data_18_15_0_lpi_1,
          buffer_bank7_data_19_15_0_lpi_1, buffer_bank7_data_20_15_0_lpi_1, buffer_bank7_data_21_15_0_lpi_1,
          buffer_bank7_data_22_15_0_lpi_1, buffer_bank7_data_23_15_0_lpi_1, buffer_bank7_data_24_15_0_lpi_1,
          buffer_bank7_data_25_15_0_lpi_1, buffer_bank7_data_26_15_0_lpi_1, buffer_bank7_data_27_15_0_lpi_1,
          buffer_bank7_data_28_15_0_lpi_1, buffer_bank7_data_29_15_0_lpi_1, buffer_bank7_data_30_15_0_lpi_1,
          buffer_bank7_data_31_15_0_lpi_1, buffer_bank7_data_32_15_0_lpi_1, buffer_bank7_data_33_15_0_lpi_1,
          buffer_bank7_data_34_15_0_lpi_1, buffer_bank7_data_35_15_0_lpi_1, buffer_bank7_data_36_15_0_lpi_1,
          buffer_bank7_data_37_15_0_lpi_1, buffer_bank7_data_38_15_0_lpi_1, buffer_bank7_data_39_15_0_lpi_1,
          buffer_bank7_data_40_15_0_lpi_1, buffer_bank7_data_41_15_0_lpi_1, buffer_bank7_data_42_15_0_lpi_1,
          buffer_bank7_data_43_15_0_lpi_1, buffer_bank7_data_44_15_0_lpi_1, buffer_bank7_data_45_15_0_lpi_1,
          buffer_bank7_data_46_15_0_lpi_1, buffer_bank7_data_47_15_0_lpi_1, buffer_bank7_data_48_15_0_lpi_1,
          buffer_bank7_data_49_15_0_lpi_1, buffer_bank7_data_50_15_0_lpi_1, buffer_bank7_data_51_15_0_lpi_1,
          buffer_bank7_data_52_15_0_lpi_1, buffer_bank7_data_53_15_0_lpi_1, buffer_bank7_data_54_15_0_lpi_1,
          buffer_bank7_data_55_15_0_lpi_1, buffer_bank7_data_56_15_0_lpi_1, buffer_bank7_data_57_15_0_lpi_1,
          buffer_bank7_data_58_15_0_lpi_1, buffer_bank7_data_59_15_0_lpi_1, buffer_bank7_data_60_15_0_lpi_1,
          buffer_bank7_data_61_15_0_lpi_1, buffer_bank7_data_62_15_0_lpi_1, (quads_in_crt_lpi_1[239:224]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_95_84 <= MUX_v_12_64_2(buffer_bank2_data_0_31_20_lpi_1,
          buffer_bank2_data_1_31_20_lpi_1, buffer_bank2_data_2_31_20_lpi_1, buffer_bank2_data_3_31_20_lpi_1,
          buffer_bank2_data_4_31_20_lpi_1, buffer_bank2_data_5_31_20_lpi_1, buffer_bank2_data_6_31_20_lpi_1,
          buffer_bank2_data_7_31_20_lpi_1, buffer_bank2_data_8_31_20_lpi_1, buffer_bank2_data_9_31_20_lpi_1,
          buffer_bank2_data_10_31_20_lpi_1, buffer_bank2_data_11_31_20_lpi_1, buffer_bank2_data_12_31_20_lpi_1,
          buffer_bank2_data_13_31_20_lpi_1, buffer_bank2_data_14_31_20_lpi_1, buffer_bank2_data_15_31_20_lpi_1,
          buffer_bank2_data_16_31_20_lpi_1, buffer_bank2_data_17_31_20_lpi_1, buffer_bank2_data_18_31_20_lpi_1,
          buffer_bank2_data_19_31_20_lpi_1, buffer_bank2_data_20_31_20_lpi_1, buffer_bank2_data_21_31_20_lpi_1,
          buffer_bank2_data_22_31_20_lpi_1, buffer_bank2_data_23_31_20_lpi_1, buffer_bank2_data_24_31_20_lpi_1,
          buffer_bank2_data_25_31_20_lpi_1, buffer_bank2_data_26_31_20_lpi_1, buffer_bank2_data_27_31_20_lpi_1,
          buffer_bank2_data_28_31_20_lpi_1, buffer_bank2_data_29_31_20_lpi_1, buffer_bank2_data_30_31_20_lpi_1,
          buffer_bank2_data_31_31_20_lpi_1, buffer_bank2_data_32_31_20_lpi_1, buffer_bank2_data_33_31_20_lpi_1,
          buffer_bank2_data_34_31_20_lpi_1, buffer_bank2_data_35_31_20_lpi_1, buffer_bank2_data_36_31_20_lpi_1,
          buffer_bank2_data_37_31_20_lpi_1, buffer_bank2_data_38_31_20_lpi_1, buffer_bank2_data_39_31_20_lpi_1,
          buffer_bank2_data_40_31_20_lpi_1, buffer_bank2_data_41_31_20_lpi_1, buffer_bank2_data_42_31_20_lpi_1,
          buffer_bank2_data_43_31_20_lpi_1, buffer_bank2_data_44_31_20_lpi_1, buffer_bank2_data_45_31_20_lpi_1,
          buffer_bank2_data_46_31_20_lpi_1, buffer_bank2_data_47_31_20_lpi_1, buffer_bank2_data_48_31_20_lpi_1,
          buffer_bank2_data_49_31_20_lpi_1, buffer_bank2_data_50_31_20_lpi_1, buffer_bank2_data_51_31_20_lpi_1,
          buffer_bank2_data_52_31_20_lpi_1, buffer_bank2_data_53_31_20_lpi_1, buffer_bank2_data_54_31_20_lpi_1,
          buffer_bank2_data_55_31_20_lpi_1, buffer_bank2_data_56_31_20_lpi_1, buffer_bank2_data_57_31_20_lpi_1,
          buffer_bank2_data_58_31_20_lpi_1, buffer_bank2_data_59_31_20_lpi_1, buffer_bank2_data_60_31_20_lpi_1,
          buffer_bank2_data_61_31_20_lpi_1, buffer_bank2_data_62_31_20_lpi_1, (quads_in_crt_lpi_1[95:84]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_223_215 <= MUX_v_9_64_2(buffer_bank6_data_0_31_23_lpi_1,
          buffer_bank6_data_1_31_23_lpi_1, buffer_bank6_data_2_31_23_lpi_1, buffer_bank6_data_3_31_23_lpi_1,
          buffer_bank6_data_4_31_23_lpi_1, buffer_bank6_data_5_31_23_lpi_1, buffer_bank6_data_6_31_23_lpi_1,
          buffer_bank6_data_7_31_23_lpi_1, buffer_bank6_data_8_31_23_lpi_1, buffer_bank6_data_9_31_23_lpi_1,
          buffer_bank6_data_10_31_23_lpi_1, buffer_bank6_data_11_31_23_lpi_1, buffer_bank6_data_12_31_23_lpi_1,
          buffer_bank6_data_13_31_23_lpi_1, buffer_bank6_data_14_31_23_lpi_1, buffer_bank6_data_15_31_23_lpi_1,
          buffer_bank6_data_16_31_23_lpi_1, buffer_bank6_data_17_31_23_lpi_1, buffer_bank6_data_18_31_23_lpi_1,
          buffer_bank6_data_19_31_23_lpi_1, buffer_bank6_data_20_31_23_lpi_1, buffer_bank6_data_21_31_23_lpi_1,
          buffer_bank6_data_22_31_23_lpi_1, buffer_bank6_data_23_31_23_lpi_1, buffer_bank6_data_24_31_23_lpi_1,
          buffer_bank6_data_25_31_23_lpi_1, buffer_bank6_data_26_31_23_lpi_1, buffer_bank6_data_27_31_23_lpi_1,
          buffer_bank6_data_28_31_23_lpi_1, buffer_bank6_data_29_31_23_lpi_1, buffer_bank6_data_30_31_23_lpi_1,
          buffer_bank6_data_31_31_23_lpi_1, buffer_bank6_data_32_31_23_lpi_1, buffer_bank6_data_33_31_23_lpi_1,
          buffer_bank6_data_34_31_23_lpi_1, buffer_bank6_data_35_31_23_lpi_1, buffer_bank6_data_36_31_23_lpi_1,
          buffer_bank6_data_37_31_23_lpi_1, buffer_bank6_data_38_31_23_lpi_1, buffer_bank6_data_39_31_23_lpi_1,
          buffer_bank6_data_40_31_23_lpi_1, buffer_bank6_data_41_31_23_lpi_1, buffer_bank6_data_42_31_23_lpi_1,
          buffer_bank6_data_43_31_23_lpi_1, buffer_bank6_data_44_31_23_lpi_1, buffer_bank6_data_45_31_23_lpi_1,
          buffer_bank6_data_46_31_23_lpi_1, buffer_bank6_data_47_31_23_lpi_1, buffer_bank6_data_48_31_23_lpi_1,
          buffer_bank6_data_49_31_23_lpi_1, buffer_bank6_data_50_31_23_lpi_1, buffer_bank6_data_51_31_23_lpi_1,
          buffer_bank6_data_52_31_23_lpi_1, buffer_bank6_data_53_31_23_lpi_1, buffer_bank6_data_54_31_23_lpi_1,
          buffer_bank6_data_55_31_23_lpi_1, buffer_bank6_data_56_31_23_lpi_1, buffer_bank6_data_57_31_23_lpi_1,
          buffer_bank6_data_58_31_23_lpi_1, buffer_bank6_data_59_31_23_lpi_1, buffer_bank6_data_60_31_23_lpi_1,
          buffer_bank6_data_61_31_23_lpi_1, buffer_bank6_data_62_31_23_lpi_1, (quads_in_crt_lpi_1[223:215]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_107_96 <= MUX_v_12_64_2(buffer_bank3_data_0_11_0_lpi_1,
          buffer_bank3_data_1_11_0_lpi_1, buffer_bank3_data_2_11_0_lpi_1, buffer_bank3_data_3_11_0_lpi_1,
          buffer_bank3_data_4_11_0_lpi_1, buffer_bank3_data_5_11_0_lpi_1, buffer_bank3_data_6_11_0_lpi_1,
          buffer_bank3_data_7_11_0_lpi_1, buffer_bank3_data_8_11_0_lpi_1, buffer_bank3_data_9_11_0_lpi_1,
          buffer_bank3_data_10_11_0_lpi_1, buffer_bank3_data_11_11_0_lpi_1, buffer_bank3_data_12_11_0_lpi_1,
          buffer_bank3_data_13_11_0_lpi_1, buffer_bank3_data_14_11_0_lpi_1, buffer_bank3_data_15_11_0_lpi_1,
          buffer_bank3_data_16_11_0_lpi_1, buffer_bank3_data_17_11_0_lpi_1, buffer_bank3_data_18_11_0_lpi_1,
          buffer_bank3_data_19_11_0_lpi_1, buffer_bank3_data_20_11_0_lpi_1, buffer_bank3_data_21_11_0_lpi_1,
          buffer_bank3_data_22_11_0_lpi_1, buffer_bank3_data_23_11_0_lpi_1, buffer_bank3_data_24_11_0_lpi_1,
          buffer_bank3_data_25_11_0_lpi_1, buffer_bank3_data_26_11_0_lpi_1, buffer_bank3_data_27_11_0_lpi_1,
          buffer_bank3_data_28_11_0_lpi_1, buffer_bank3_data_29_11_0_lpi_1, buffer_bank3_data_30_11_0_lpi_1,
          buffer_bank3_data_31_11_0_lpi_1, buffer_bank3_data_32_11_0_lpi_1, buffer_bank3_data_33_11_0_lpi_1,
          buffer_bank3_data_34_11_0_lpi_1, buffer_bank3_data_35_11_0_lpi_1, buffer_bank3_data_36_11_0_lpi_1,
          buffer_bank3_data_37_11_0_lpi_1, buffer_bank3_data_38_11_0_lpi_1, buffer_bank3_data_39_11_0_lpi_1,
          buffer_bank3_data_40_11_0_lpi_1, buffer_bank3_data_41_11_0_lpi_1, buffer_bank3_data_42_11_0_lpi_1,
          buffer_bank3_data_43_11_0_lpi_1, buffer_bank3_data_44_11_0_lpi_1, buffer_bank3_data_45_11_0_lpi_1,
          buffer_bank3_data_46_11_0_lpi_1, buffer_bank3_data_47_11_0_lpi_1, buffer_bank3_data_48_11_0_lpi_1,
          buffer_bank3_data_49_11_0_lpi_1, buffer_bank3_data_50_11_0_lpi_1, buffer_bank3_data_51_11_0_lpi_1,
          buffer_bank3_data_52_11_0_lpi_1, buffer_bank3_data_53_11_0_lpi_1, buffer_bank3_data_54_11_0_lpi_1,
          buffer_bank3_data_55_11_0_lpi_1, buffer_bank3_data_56_11_0_lpi_1, buffer_bank3_data_57_11_0_lpi_1,
          buffer_bank3_data_58_11_0_lpi_1, buffer_bank3_data_59_11_0_lpi_1, buffer_bank3_data_60_11_0_lpi_1,
          buffer_bank3_data_61_11_0_lpi_1, buffer_bank3_data_62_11_0_lpi_1, (quads_in_crt_lpi_1[107:96]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_214_192 <= MUX_v_23_64_2(buffer_bank6_data_0_22_0_lpi_1,
          buffer_bank6_data_1_22_0_lpi_1, buffer_bank6_data_2_22_0_lpi_1, buffer_bank6_data_3_22_0_lpi_1,
          buffer_bank6_data_4_22_0_lpi_1, buffer_bank6_data_5_22_0_lpi_1, buffer_bank6_data_6_22_0_lpi_1,
          buffer_bank6_data_7_22_0_lpi_1, buffer_bank6_data_8_22_0_lpi_1, buffer_bank6_data_9_22_0_lpi_1,
          buffer_bank6_data_10_22_0_lpi_1, buffer_bank6_data_11_22_0_lpi_1, buffer_bank6_data_12_22_0_lpi_1,
          buffer_bank6_data_13_22_0_lpi_1, buffer_bank6_data_14_22_0_lpi_1, buffer_bank6_data_15_22_0_lpi_1,
          buffer_bank6_data_16_22_0_lpi_1, buffer_bank6_data_17_22_0_lpi_1, buffer_bank6_data_18_22_0_lpi_1,
          buffer_bank6_data_19_22_0_lpi_1, buffer_bank6_data_20_22_0_lpi_1, buffer_bank6_data_21_22_0_lpi_1,
          buffer_bank6_data_22_22_0_lpi_1, buffer_bank6_data_23_22_0_lpi_1, buffer_bank6_data_24_22_0_lpi_1,
          buffer_bank6_data_25_22_0_lpi_1, buffer_bank6_data_26_22_0_lpi_1, buffer_bank6_data_27_22_0_lpi_1,
          buffer_bank6_data_28_22_0_lpi_1, buffer_bank6_data_29_22_0_lpi_1, buffer_bank6_data_30_22_0_lpi_1,
          buffer_bank6_data_31_22_0_lpi_1, buffer_bank6_data_32_22_0_lpi_1, buffer_bank6_data_33_22_0_lpi_1,
          buffer_bank6_data_34_22_0_lpi_1, buffer_bank6_data_35_22_0_lpi_1, buffer_bank6_data_36_22_0_lpi_1,
          buffer_bank6_data_37_22_0_lpi_1, buffer_bank6_data_38_22_0_lpi_1, buffer_bank6_data_39_22_0_lpi_1,
          buffer_bank6_data_40_22_0_lpi_1, buffer_bank6_data_41_22_0_lpi_1, buffer_bank6_data_42_22_0_lpi_1,
          buffer_bank6_data_43_22_0_lpi_1, buffer_bank6_data_44_22_0_lpi_1, buffer_bank6_data_45_22_0_lpi_1,
          buffer_bank6_data_46_22_0_lpi_1, buffer_bank6_data_47_22_0_lpi_1, buffer_bank6_data_48_22_0_lpi_1,
          buffer_bank6_data_49_22_0_lpi_1, buffer_bank6_data_50_22_0_lpi_1, buffer_bank6_data_51_22_0_lpi_1,
          buffer_bank6_data_52_22_0_lpi_1, buffer_bank6_data_53_22_0_lpi_1, buffer_bank6_data_54_22_0_lpi_1,
          buffer_bank6_data_55_22_0_lpi_1, buffer_bank6_data_56_22_0_lpi_1, buffer_bank6_data_57_22_0_lpi_1,
          buffer_bank6_data_58_22_0_lpi_1, buffer_bank6_data_59_22_0_lpi_1, buffer_bank6_data_60_22_0_lpi_1,
          buffer_bank6_data_61_22_0_lpi_1, buffer_bank6_data_62_22_0_lpi_1, (quads_in_crt_lpi_1[214:192]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_110_108 <= MUX_v_3_64_2(buffer_bank3_data_0_14_12_lpi_1,
          buffer_bank3_data_1_14_12_lpi_1, buffer_bank3_data_2_14_12_lpi_1, buffer_bank3_data_3_14_12_lpi_1,
          buffer_bank3_data_4_14_12_lpi_1, buffer_bank3_data_5_14_12_lpi_1, buffer_bank3_data_6_14_12_lpi_1,
          buffer_bank3_data_7_14_12_lpi_1, buffer_bank3_data_8_14_12_lpi_1, buffer_bank3_data_9_14_12_lpi_1,
          buffer_bank3_data_10_14_12_lpi_1, buffer_bank3_data_11_14_12_lpi_1, buffer_bank3_data_12_14_12_lpi_1,
          buffer_bank3_data_13_14_12_lpi_1, buffer_bank3_data_14_14_12_lpi_1, buffer_bank3_data_15_14_12_lpi_1,
          buffer_bank3_data_16_14_12_lpi_1, buffer_bank3_data_17_14_12_lpi_1, buffer_bank3_data_18_14_12_lpi_1,
          buffer_bank3_data_19_14_12_lpi_1, buffer_bank3_data_20_14_12_lpi_1, buffer_bank3_data_21_14_12_lpi_1,
          buffer_bank3_data_22_14_12_lpi_1, buffer_bank3_data_23_14_12_lpi_1, buffer_bank3_data_24_14_12_lpi_1,
          buffer_bank3_data_25_14_12_lpi_1, buffer_bank3_data_26_14_12_lpi_1, buffer_bank3_data_27_14_12_lpi_1,
          buffer_bank3_data_28_14_12_lpi_1, buffer_bank3_data_29_14_12_lpi_1, buffer_bank3_data_30_14_12_lpi_1,
          buffer_bank3_data_31_14_12_lpi_1, buffer_bank3_data_32_14_12_lpi_1, buffer_bank3_data_33_14_12_lpi_1,
          buffer_bank3_data_34_14_12_lpi_1, buffer_bank3_data_35_14_12_lpi_1, buffer_bank3_data_36_14_12_lpi_1,
          buffer_bank3_data_37_14_12_lpi_1, buffer_bank3_data_38_14_12_lpi_1, buffer_bank3_data_39_14_12_lpi_1,
          buffer_bank3_data_40_14_12_lpi_1, buffer_bank3_data_41_14_12_lpi_1, buffer_bank3_data_42_14_12_lpi_1,
          buffer_bank3_data_43_14_12_lpi_1, buffer_bank3_data_44_14_12_lpi_1, buffer_bank3_data_45_14_12_lpi_1,
          buffer_bank3_data_46_14_12_lpi_1, buffer_bank3_data_47_14_12_lpi_1, buffer_bank3_data_48_14_12_lpi_1,
          buffer_bank3_data_49_14_12_lpi_1, buffer_bank3_data_50_14_12_lpi_1, buffer_bank3_data_51_14_12_lpi_1,
          buffer_bank3_data_52_14_12_lpi_1, buffer_bank3_data_53_14_12_lpi_1, buffer_bank3_data_54_14_12_lpi_1,
          buffer_bank3_data_55_14_12_lpi_1, buffer_bank3_data_56_14_12_lpi_1, buffer_bank3_data_57_14_12_lpi_1,
          buffer_bank3_data_58_14_12_lpi_1, buffer_bank3_data_59_14_12_lpi_1, buffer_bank3_data_60_14_12_lpi_1,
          buffer_bank3_data_61_14_12_lpi_1, buffer_bank3_data_62_14_12_lpi_1, (quads_in_crt_lpi_1[110:108]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_191_190 <= MUX_v_2_64_2(buffer_bank5_data_0_31_30_lpi_1,
          buffer_bank5_data_1_31_30_lpi_1, buffer_bank5_data_2_31_30_lpi_1, buffer_bank5_data_3_31_30_lpi_1,
          buffer_bank5_data_4_31_30_lpi_1, buffer_bank5_data_5_31_30_lpi_1, buffer_bank5_data_6_31_30_lpi_1,
          buffer_bank5_data_7_31_30_lpi_1, buffer_bank5_data_8_31_30_lpi_1, buffer_bank5_data_9_31_30_lpi_1,
          buffer_bank5_data_10_31_30_lpi_1, buffer_bank5_data_11_31_30_lpi_1, buffer_bank5_data_12_31_30_lpi_1,
          buffer_bank5_data_13_31_30_lpi_1, buffer_bank5_data_14_31_30_lpi_1, buffer_bank5_data_15_31_30_lpi_1,
          buffer_bank5_data_16_31_30_lpi_1, buffer_bank5_data_17_31_30_lpi_1, buffer_bank5_data_18_31_30_lpi_1,
          buffer_bank5_data_19_31_30_lpi_1, buffer_bank5_data_20_31_30_lpi_1, buffer_bank5_data_21_31_30_lpi_1,
          buffer_bank5_data_22_31_30_lpi_1, buffer_bank5_data_23_31_30_lpi_1, buffer_bank5_data_24_31_30_lpi_1,
          buffer_bank5_data_25_31_30_lpi_1, buffer_bank5_data_26_31_30_lpi_1, buffer_bank5_data_27_31_30_lpi_1,
          buffer_bank5_data_28_31_30_lpi_1, buffer_bank5_data_29_31_30_lpi_1, buffer_bank5_data_30_31_30_lpi_1,
          buffer_bank5_data_31_31_30_lpi_1, buffer_bank5_data_32_31_30_lpi_1, buffer_bank5_data_33_31_30_lpi_1,
          buffer_bank5_data_34_31_30_lpi_1, buffer_bank5_data_35_31_30_lpi_1, buffer_bank5_data_36_31_30_lpi_1,
          buffer_bank5_data_37_31_30_lpi_1, buffer_bank5_data_38_31_30_lpi_1, buffer_bank5_data_39_31_30_lpi_1,
          buffer_bank5_data_40_31_30_lpi_1, buffer_bank5_data_41_31_30_lpi_1, buffer_bank5_data_42_31_30_lpi_1,
          buffer_bank5_data_43_31_30_lpi_1, buffer_bank5_data_44_31_30_lpi_1, buffer_bank5_data_45_31_30_lpi_1,
          buffer_bank5_data_46_31_30_lpi_1, buffer_bank5_data_47_31_30_lpi_1, buffer_bank5_data_48_31_30_lpi_1,
          buffer_bank5_data_49_31_30_lpi_1, buffer_bank5_data_50_31_30_lpi_1, buffer_bank5_data_51_31_30_lpi_1,
          buffer_bank5_data_52_31_30_lpi_1, buffer_bank5_data_53_31_30_lpi_1, buffer_bank5_data_54_31_30_lpi_1,
          buffer_bank5_data_55_31_30_lpi_1, buffer_bank5_data_56_31_30_lpi_1, buffer_bank5_data_57_31_30_lpi_1,
          buffer_bank5_data_58_31_30_lpi_1, buffer_bank5_data_59_31_30_lpi_1, buffer_bank5_data_60_31_30_lpi_1,
          buffer_bank5_data_61_31_30_lpi_1, buffer_bank5_data_62_31_30_lpi_1, (quads_in_crt_lpi_1[191:190]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_111 <= MUX_s_1_64_2(buffer_bank3_data_0_15_lpi_1, buffer_bank3_data_1_15_lpi_1,
          buffer_bank3_data_2_15_lpi_1, buffer_bank3_data_3_15_lpi_1, buffer_bank3_data_4_15_lpi_1,
          buffer_bank3_data_5_15_lpi_1, buffer_bank3_data_6_15_lpi_1, buffer_bank3_data_7_15_lpi_1,
          buffer_bank3_data_8_15_lpi_1, buffer_bank3_data_9_15_lpi_1, buffer_bank3_data_10_15_lpi_1,
          buffer_bank3_data_11_15_lpi_1, buffer_bank3_data_12_15_lpi_1, buffer_bank3_data_13_15_lpi_1,
          buffer_bank3_data_14_15_lpi_1, buffer_bank3_data_15_15_lpi_1, buffer_bank3_data_16_15_lpi_1,
          buffer_bank3_data_17_15_lpi_1, buffer_bank3_data_18_15_lpi_1, buffer_bank3_data_19_15_lpi_1,
          buffer_bank3_data_20_15_lpi_1, buffer_bank3_data_21_15_lpi_1, buffer_bank3_data_22_15_lpi_1,
          buffer_bank3_data_23_15_lpi_1, buffer_bank3_data_24_15_lpi_1, buffer_bank3_data_25_15_lpi_1,
          buffer_bank3_data_26_15_lpi_1, buffer_bank3_data_27_15_lpi_1, buffer_bank3_data_28_15_lpi_1,
          buffer_bank3_data_29_15_lpi_1, buffer_bank3_data_30_15_lpi_1, buffer_bank3_data_31_15_lpi_1,
          buffer_bank3_data_32_15_lpi_1, buffer_bank3_data_33_15_lpi_1, buffer_bank3_data_34_15_lpi_1,
          buffer_bank3_data_35_15_lpi_1, buffer_bank3_data_36_15_lpi_1, buffer_bank3_data_37_15_lpi_1,
          buffer_bank3_data_38_15_lpi_1, buffer_bank3_data_39_15_lpi_1, buffer_bank3_data_40_15_lpi_1,
          buffer_bank3_data_41_15_lpi_1, buffer_bank3_data_42_15_lpi_1, buffer_bank3_data_43_15_lpi_1,
          buffer_bank3_data_44_15_lpi_1, buffer_bank3_data_45_15_lpi_1, buffer_bank3_data_46_15_lpi_1,
          buffer_bank3_data_47_15_lpi_1, buffer_bank3_data_48_15_lpi_1, buffer_bank3_data_49_15_lpi_1,
          buffer_bank3_data_50_15_lpi_1, buffer_bank3_data_51_15_lpi_1, buffer_bank3_data_52_15_lpi_1,
          buffer_bank3_data_53_15_lpi_1, buffer_bank3_data_54_15_lpi_1, buffer_bank3_data_55_15_lpi_1,
          buffer_bank3_data_56_15_lpi_1, buffer_bank3_data_57_15_lpi_1, buffer_bank3_data_58_15_lpi_1,
          buffer_bank3_data_59_15_lpi_1, buffer_bank3_data_60_15_lpi_1, buffer_bank3_data_61_15_lpi_1,
          buffer_bank3_data_62_15_lpi_1, (quads_in_crt_lpi_1[111]), for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_189_164 <= MUX_v_26_64_2(buffer_bank5_data_0_29_4_lpi_1,
          buffer_bank5_data_1_29_4_lpi_1, buffer_bank5_data_2_29_4_lpi_1, buffer_bank5_data_3_29_4_lpi_1,
          buffer_bank5_data_4_29_4_lpi_1, buffer_bank5_data_5_29_4_lpi_1, buffer_bank5_data_6_29_4_lpi_1,
          buffer_bank5_data_7_29_4_lpi_1, buffer_bank5_data_8_29_4_lpi_1, buffer_bank5_data_9_29_4_lpi_1,
          buffer_bank5_data_10_29_4_lpi_1, buffer_bank5_data_11_29_4_lpi_1, buffer_bank5_data_12_29_4_lpi_1,
          buffer_bank5_data_13_29_4_lpi_1, buffer_bank5_data_14_29_4_lpi_1, buffer_bank5_data_15_29_4_lpi_1,
          buffer_bank5_data_16_29_4_lpi_1, buffer_bank5_data_17_29_4_lpi_1, buffer_bank5_data_18_29_4_lpi_1,
          buffer_bank5_data_19_29_4_lpi_1, buffer_bank5_data_20_29_4_lpi_1, buffer_bank5_data_21_29_4_lpi_1,
          buffer_bank5_data_22_29_4_lpi_1, buffer_bank5_data_23_29_4_lpi_1, buffer_bank5_data_24_29_4_lpi_1,
          buffer_bank5_data_25_29_4_lpi_1, buffer_bank5_data_26_29_4_lpi_1, buffer_bank5_data_27_29_4_lpi_1,
          buffer_bank5_data_28_29_4_lpi_1, buffer_bank5_data_29_29_4_lpi_1, buffer_bank5_data_30_29_4_lpi_1,
          buffer_bank5_data_31_29_4_lpi_1, buffer_bank5_data_32_29_4_lpi_1, buffer_bank5_data_33_29_4_lpi_1,
          buffer_bank5_data_34_29_4_lpi_1, buffer_bank5_data_35_29_4_lpi_1, buffer_bank5_data_36_29_4_lpi_1,
          buffer_bank5_data_37_29_4_lpi_1, buffer_bank5_data_38_29_4_lpi_1, buffer_bank5_data_39_29_4_lpi_1,
          buffer_bank5_data_40_29_4_lpi_1, buffer_bank5_data_41_29_4_lpi_1, buffer_bank5_data_42_29_4_lpi_1,
          buffer_bank5_data_43_29_4_lpi_1, buffer_bank5_data_44_29_4_lpi_1, buffer_bank5_data_45_29_4_lpi_1,
          buffer_bank5_data_46_29_4_lpi_1, buffer_bank5_data_47_29_4_lpi_1, buffer_bank5_data_48_29_4_lpi_1,
          buffer_bank5_data_49_29_4_lpi_1, buffer_bank5_data_50_29_4_lpi_1, buffer_bank5_data_51_29_4_lpi_1,
          buffer_bank5_data_52_29_4_lpi_1, buffer_bank5_data_53_29_4_lpi_1, buffer_bank5_data_54_29_4_lpi_1,
          buffer_bank5_data_55_29_4_lpi_1, buffer_bank5_data_56_29_4_lpi_1, buffer_bank5_data_57_29_4_lpi_1,
          buffer_bank5_data_58_29_4_lpi_1, buffer_bank5_data_59_29_4_lpi_1, buffer_bank5_data_60_29_4_lpi_1,
          buffer_bank5_data_61_29_4_lpi_1, buffer_bank5_data_62_29_4_lpi_1, (quads_in_crt_lpi_1[189:164]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_127_112 <= MUX_v_16_64_2(buffer_bank3_data_0_31_16_lpi_1,
          buffer_bank3_data_1_31_16_lpi_1, buffer_bank3_data_2_31_16_lpi_1, buffer_bank3_data_3_31_16_lpi_1,
          buffer_bank3_data_4_31_16_lpi_1, buffer_bank3_data_5_31_16_lpi_1, buffer_bank3_data_6_31_16_lpi_1,
          buffer_bank3_data_7_31_16_lpi_1, buffer_bank3_data_8_31_16_lpi_1, buffer_bank3_data_9_31_16_lpi_1,
          buffer_bank3_data_10_31_16_lpi_1, buffer_bank3_data_11_31_16_lpi_1, buffer_bank3_data_12_31_16_lpi_1,
          buffer_bank3_data_13_31_16_lpi_1, buffer_bank3_data_14_31_16_lpi_1, buffer_bank3_data_15_31_16_lpi_1,
          buffer_bank3_data_16_31_16_lpi_1, buffer_bank3_data_17_31_16_lpi_1, buffer_bank3_data_18_31_16_lpi_1,
          buffer_bank3_data_19_31_16_lpi_1, buffer_bank3_data_20_31_16_lpi_1, buffer_bank3_data_21_31_16_lpi_1,
          buffer_bank3_data_22_31_16_lpi_1, buffer_bank3_data_23_31_16_lpi_1, buffer_bank3_data_24_31_16_lpi_1,
          buffer_bank3_data_25_31_16_lpi_1, buffer_bank3_data_26_31_16_lpi_1, buffer_bank3_data_27_31_16_lpi_1,
          buffer_bank3_data_28_31_16_lpi_1, buffer_bank3_data_29_31_16_lpi_1, buffer_bank3_data_30_31_16_lpi_1,
          buffer_bank3_data_31_31_16_lpi_1, buffer_bank3_data_32_31_16_lpi_1, buffer_bank3_data_33_31_16_lpi_1,
          buffer_bank3_data_34_31_16_lpi_1, buffer_bank3_data_35_31_16_lpi_1, buffer_bank3_data_36_31_16_lpi_1,
          buffer_bank3_data_37_31_16_lpi_1, buffer_bank3_data_38_31_16_lpi_1, buffer_bank3_data_39_31_16_lpi_1,
          buffer_bank3_data_40_31_16_lpi_1, buffer_bank3_data_41_31_16_lpi_1, buffer_bank3_data_42_31_16_lpi_1,
          buffer_bank3_data_43_31_16_lpi_1, buffer_bank3_data_44_31_16_lpi_1, buffer_bank3_data_45_31_16_lpi_1,
          buffer_bank3_data_46_31_16_lpi_1, buffer_bank3_data_47_31_16_lpi_1, buffer_bank3_data_48_31_16_lpi_1,
          buffer_bank3_data_49_31_16_lpi_1, buffer_bank3_data_50_31_16_lpi_1, buffer_bank3_data_51_31_16_lpi_1,
          buffer_bank3_data_52_31_16_lpi_1, buffer_bank3_data_53_31_16_lpi_1, buffer_bank3_data_54_31_16_lpi_1,
          buffer_bank3_data_55_31_16_lpi_1, buffer_bank3_data_56_31_16_lpi_1, buffer_bank3_data_57_31_16_lpi_1,
          buffer_bank3_data_58_31_16_lpi_1, buffer_bank3_data_59_31_16_lpi_1, buffer_bank3_data_60_31_16_lpi_1,
          buffer_bank3_data_61_31_16_lpi_1, buffer_bank3_data_62_31_16_lpi_1, (quads_in_crt_lpi_1[127:112]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_163_160 <= MUX_v_4_64_2(buffer_bank5_data_0_3_0_lpi_1,
          buffer_bank5_data_1_3_0_lpi_1, buffer_bank5_data_2_3_0_lpi_1, buffer_bank5_data_3_3_0_lpi_1,
          buffer_bank5_data_4_3_0_lpi_1, buffer_bank5_data_5_3_0_lpi_1, buffer_bank5_data_6_3_0_lpi_1,
          buffer_bank5_data_7_3_0_lpi_1, buffer_bank5_data_8_3_0_lpi_1, buffer_bank5_data_9_3_0_lpi_1,
          buffer_bank5_data_10_3_0_lpi_1, buffer_bank5_data_11_3_0_lpi_1, buffer_bank5_data_12_3_0_lpi_1,
          buffer_bank5_data_13_3_0_lpi_1, buffer_bank5_data_14_3_0_lpi_1, buffer_bank5_data_15_3_0_lpi_1,
          buffer_bank5_data_16_3_0_lpi_1, buffer_bank5_data_17_3_0_lpi_1, buffer_bank5_data_18_3_0_lpi_1,
          buffer_bank5_data_19_3_0_lpi_1, buffer_bank5_data_20_3_0_lpi_1, buffer_bank5_data_21_3_0_lpi_1,
          buffer_bank5_data_22_3_0_lpi_1, buffer_bank5_data_23_3_0_lpi_1, buffer_bank5_data_24_3_0_lpi_1,
          buffer_bank5_data_25_3_0_lpi_1, buffer_bank5_data_26_3_0_lpi_1, buffer_bank5_data_27_3_0_lpi_1,
          buffer_bank5_data_28_3_0_lpi_1, buffer_bank5_data_29_3_0_lpi_1, buffer_bank5_data_30_3_0_lpi_1,
          buffer_bank5_data_31_3_0_lpi_1, buffer_bank5_data_32_3_0_lpi_1, buffer_bank5_data_33_3_0_lpi_1,
          buffer_bank5_data_34_3_0_lpi_1, buffer_bank5_data_35_3_0_lpi_1, buffer_bank5_data_36_3_0_lpi_1,
          buffer_bank5_data_37_3_0_lpi_1, buffer_bank5_data_38_3_0_lpi_1, buffer_bank5_data_39_3_0_lpi_1,
          buffer_bank5_data_40_3_0_lpi_1, buffer_bank5_data_41_3_0_lpi_1, buffer_bank5_data_42_3_0_lpi_1,
          buffer_bank5_data_43_3_0_lpi_1, buffer_bank5_data_44_3_0_lpi_1, buffer_bank5_data_45_3_0_lpi_1,
          buffer_bank5_data_46_3_0_lpi_1, buffer_bank5_data_47_3_0_lpi_1, buffer_bank5_data_48_3_0_lpi_1,
          buffer_bank5_data_49_3_0_lpi_1, buffer_bank5_data_50_3_0_lpi_1, buffer_bank5_data_51_3_0_lpi_1,
          buffer_bank5_data_52_3_0_lpi_1, buffer_bank5_data_53_3_0_lpi_1, buffer_bank5_data_54_3_0_lpi_1,
          buffer_bank5_data_55_3_0_lpi_1, buffer_bank5_data_56_3_0_lpi_1, buffer_bank5_data_57_3_0_lpi_1,
          buffer_bank5_data_58_3_0_lpi_1, buffer_bank5_data_59_3_0_lpi_1, buffer_bank5_data_60_3_0_lpi_1,
          buffer_bank5_data_61_3_0_lpi_1, buffer_bank5_data_62_3_0_lpi_1, (quads_in_crt_lpi_1[163:160]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_137_128 <= MUX_v_10_64_2(buffer_bank4_data_0_9_0_lpi_1,
          buffer_bank4_data_1_9_0_lpi_1, buffer_bank4_data_2_9_0_lpi_1, buffer_bank4_data_3_9_0_lpi_1,
          buffer_bank4_data_4_9_0_lpi_1, buffer_bank4_data_5_9_0_lpi_1, buffer_bank4_data_6_9_0_lpi_1,
          buffer_bank4_data_7_9_0_lpi_1, buffer_bank4_data_8_9_0_lpi_1, buffer_bank4_data_9_9_0_lpi_1,
          buffer_bank4_data_10_9_0_lpi_1, buffer_bank4_data_11_9_0_lpi_1, buffer_bank4_data_12_9_0_lpi_1,
          buffer_bank4_data_13_9_0_lpi_1, buffer_bank4_data_14_9_0_lpi_1, buffer_bank4_data_15_9_0_lpi_1,
          buffer_bank4_data_16_9_0_lpi_1, buffer_bank4_data_17_9_0_lpi_1, buffer_bank4_data_18_9_0_lpi_1,
          buffer_bank4_data_19_9_0_lpi_1, buffer_bank4_data_20_9_0_lpi_1, buffer_bank4_data_21_9_0_lpi_1,
          buffer_bank4_data_22_9_0_lpi_1, buffer_bank4_data_23_9_0_lpi_1, buffer_bank4_data_24_9_0_lpi_1,
          buffer_bank4_data_25_9_0_lpi_1, buffer_bank4_data_26_9_0_lpi_1, buffer_bank4_data_27_9_0_lpi_1,
          buffer_bank4_data_28_9_0_lpi_1, buffer_bank4_data_29_9_0_lpi_1, buffer_bank4_data_30_9_0_lpi_1,
          buffer_bank4_data_31_9_0_lpi_1, buffer_bank4_data_32_9_0_lpi_1, buffer_bank4_data_33_9_0_lpi_1,
          buffer_bank4_data_34_9_0_lpi_1, buffer_bank4_data_35_9_0_lpi_1, buffer_bank4_data_36_9_0_lpi_1,
          buffer_bank4_data_37_9_0_lpi_1, buffer_bank4_data_38_9_0_lpi_1, buffer_bank4_data_39_9_0_lpi_1,
          buffer_bank4_data_40_9_0_lpi_1, buffer_bank4_data_41_9_0_lpi_1, buffer_bank4_data_42_9_0_lpi_1,
          buffer_bank4_data_43_9_0_lpi_1, buffer_bank4_data_44_9_0_lpi_1, buffer_bank4_data_45_9_0_lpi_1,
          buffer_bank4_data_46_9_0_lpi_1, buffer_bank4_data_47_9_0_lpi_1, buffer_bank4_data_48_9_0_lpi_1,
          buffer_bank4_data_49_9_0_lpi_1, buffer_bank4_data_50_9_0_lpi_1, buffer_bank4_data_51_9_0_lpi_1,
          buffer_bank4_data_52_9_0_lpi_1, buffer_bank4_data_53_9_0_lpi_1, buffer_bank4_data_54_9_0_lpi_1,
          buffer_bank4_data_55_9_0_lpi_1, buffer_bank4_data_56_9_0_lpi_1, buffer_bank4_data_57_9_0_lpi_1,
          buffer_bank4_data_58_9_0_lpi_1, buffer_bank4_data_59_9_0_lpi_1, buffer_bank4_data_60_9_0_lpi_1,
          buffer_bank4_data_61_9_0_lpi_1, buffer_bank4_data_62_9_0_lpi_1, (quads_in_crt_lpi_1[137:128]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
      quads_out_rsci_idat_159_138 <= MUX_v_22_64_2(buffer_bank4_data_0_31_10_lpi_1,
          buffer_bank4_data_1_31_10_lpi_1, buffer_bank4_data_2_31_10_lpi_1, buffer_bank4_data_3_31_10_lpi_1,
          buffer_bank4_data_4_31_10_lpi_1, buffer_bank4_data_5_31_10_lpi_1, buffer_bank4_data_6_31_10_lpi_1,
          buffer_bank4_data_7_31_10_lpi_1, buffer_bank4_data_8_31_10_lpi_1, buffer_bank4_data_9_31_10_lpi_1,
          buffer_bank4_data_10_31_10_lpi_1, buffer_bank4_data_11_31_10_lpi_1, buffer_bank4_data_12_31_10_lpi_1,
          buffer_bank4_data_13_31_10_lpi_1, buffer_bank4_data_14_31_10_lpi_1, buffer_bank4_data_15_31_10_lpi_1,
          buffer_bank4_data_16_31_10_lpi_1, buffer_bank4_data_17_31_10_lpi_1, buffer_bank4_data_18_31_10_lpi_1,
          buffer_bank4_data_19_31_10_lpi_1, buffer_bank4_data_20_31_10_lpi_1, buffer_bank4_data_21_31_10_lpi_1,
          buffer_bank4_data_22_31_10_lpi_1, buffer_bank4_data_23_31_10_lpi_1, buffer_bank4_data_24_31_10_lpi_1,
          buffer_bank4_data_25_31_10_lpi_1, buffer_bank4_data_26_31_10_lpi_1, buffer_bank4_data_27_31_10_lpi_1,
          buffer_bank4_data_28_31_10_lpi_1, buffer_bank4_data_29_31_10_lpi_1, buffer_bank4_data_30_31_10_lpi_1,
          buffer_bank4_data_31_31_10_lpi_1, buffer_bank4_data_32_31_10_lpi_1, buffer_bank4_data_33_31_10_lpi_1,
          buffer_bank4_data_34_31_10_lpi_1, buffer_bank4_data_35_31_10_lpi_1, buffer_bank4_data_36_31_10_lpi_1,
          buffer_bank4_data_37_31_10_lpi_1, buffer_bank4_data_38_31_10_lpi_1, buffer_bank4_data_39_31_10_lpi_1,
          buffer_bank4_data_40_31_10_lpi_1, buffer_bank4_data_41_31_10_lpi_1, buffer_bank4_data_42_31_10_lpi_1,
          buffer_bank4_data_43_31_10_lpi_1, buffer_bank4_data_44_31_10_lpi_1, buffer_bank4_data_45_31_10_lpi_1,
          buffer_bank4_data_46_31_10_lpi_1, buffer_bank4_data_47_31_10_lpi_1, buffer_bank4_data_48_31_10_lpi_1,
          buffer_bank4_data_49_31_10_lpi_1, buffer_bank4_data_50_31_10_lpi_1, buffer_bank4_data_51_31_10_lpi_1,
          buffer_bank4_data_52_31_10_lpi_1, buffer_bank4_data_53_31_10_lpi_1, buffer_bank4_data_54_31_10_lpi_1,
          buffer_bank4_data_55_31_10_lpi_1, buffer_bank4_data_56_31_10_lpi_1, buffer_bank4_data_57_31_10_lpi_1,
          buffer_bank4_data_58_31_10_lpi_1, buffer_bank4_data_59_31_10_lpi_1, buffer_bank4_data_60_31_10_lpi_1,
          buffer_bank4_data_61_31_10_lpi_1, buffer_bank4_data_62_31_10_lpi_1, (quads_in_crt_lpi_1[159:138]),
          for_1_for_quad_idx_lpi_1_dfm_5_0_1);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exit_for_1_sva <= 1'b1;
      sfi_exit_for_1_lpi_1 <= 1'b0;
    end
    else if ( for_1_and_1901_cse ) begin
      exitL_exit_for_1_sva <= mux_89_cse;
      sfi_exit_for_1_lpi_1 <= sfi_exit_for_1_lpi_1 & (~ for_1_for_1_and_1_tmp);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_lpi_1_dfm_12_0 <= 13'b0000000000000;
    end
    else if ( run_wen & or_1_cse & main_stage_0_2 & exitL_exit_for_1_sva ) begin
      paramsIn_crt_lpi_1_dfm_12_0 <= paramsIn_rsci_idat_mxwt[12:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_i_6_0_lpi_1_dfm_1_5_0 <= 6'b000000;
    end
    else if ( (~ (mux_93_nl)) & run_wen ) begin
      for_i_6_0_lpi_1_dfm_1_5_0 <= MUX_v_6_2_2(6'b000000, (for_acc_1_tmp[5:0]), (for_1_not_3868_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_for_sva <= 1'b0;
      quads_in_crt_lpi_1 <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( for_and_123_cse ) begin
      exit_for_sva <= operator_33_true_operator_33_true_and_tmp;
      quads_in_crt_lpi_1 <= quads_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exit_for_1_lpi_1_dfm_1 <= 2'b00;
    end
    else if ( (mux_97_nl) & run_wen ) begin
      lfst_exit_for_1_lpi_1_dfm_1 <= for_1_for_1_and_4_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_1_read_request_lpi_1 <= 43'b0000000000000000000000000000000000000000000;
    end
    else if ( (mux_106_nl) & for_1_and_1901_cse ) begin
      for_1_read_request_lpi_1 <= MUX_v_43_2_2((for_for_and_nl), z_out, for_1_and_1900_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_0_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_0_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_0_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_0_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_0_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_0_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_0_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_0_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_0_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_0_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_0_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_0_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_0_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_0_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_0_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_0_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_0_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_0_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_0_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_0_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_0_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_0_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_0_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_0_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_0_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_0_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_0_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_0_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_0_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_0_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_cse ) begin
      buffer_bank11_data_0_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_0_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_0_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_0_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_0_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_0_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_0_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_0_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_0_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_0_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_0_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_0_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_0_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_0_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_0_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_0_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_0_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_0_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_0_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_0_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_0_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_0_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_0_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_0_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_0_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_0_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_0_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_0_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_0_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_0_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_1_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_1_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_1_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_1_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_1_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_1_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_1_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_1_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_1_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_1_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_1_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_1_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_1_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_1_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_1_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_1_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_1_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_1_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_1_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_1_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_1_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_1_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_1_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_1_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_1_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_1_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_1_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_1_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_1_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_1_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_1_cse ) begin
      buffer_bank11_data_1_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_1_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_1_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_1_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_1_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_1_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_1_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_1_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_1_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_1_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_1_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_1_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_1_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_1_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_1_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_1_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_1_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_1_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_1_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_1_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_1_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_1_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_1_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_1_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_1_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_1_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_1_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_1_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_1_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_1_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_2_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_2_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_2_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_2_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_2_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_2_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_2_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_2_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_2_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_2_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_2_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_2_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_2_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_2_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_2_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_2_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_2_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_2_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_2_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_2_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_2_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_2_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_2_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_2_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_2_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_2_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_2_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_2_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_2_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_2_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_2_cse ) begin
      buffer_bank11_data_2_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_2_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_2_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_2_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_2_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_2_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_2_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_2_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_2_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_2_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_2_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_2_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_2_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_2_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_2_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_2_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_2_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_2_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_2_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_2_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_2_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_2_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_2_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_2_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_2_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_2_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_2_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_2_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_2_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_2_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_3_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_3_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_3_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_3_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_3_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_3_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_3_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_3_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_3_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_3_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_3_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_3_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_3_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_3_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_3_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_3_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_3_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_3_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_3_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_3_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_3_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_3_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_3_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_3_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_3_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_3_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_3_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_3_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_3_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_3_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_3_cse ) begin
      buffer_bank11_data_3_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_3_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_3_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_3_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_3_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_3_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_3_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_3_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_3_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_3_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_3_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_3_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_3_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_3_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_3_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_3_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_3_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_3_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_3_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_3_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_3_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_3_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_3_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_3_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_3_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_3_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_3_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_3_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_3_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_3_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_4_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_4_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_4_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_4_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_4_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_4_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_4_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_4_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_4_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_4_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_4_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_4_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_4_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_4_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_4_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_4_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_4_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_4_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_4_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_4_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_4_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_4_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_4_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_4_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_4_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_4_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_4_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_4_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_4_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_4_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_4_cse ) begin
      buffer_bank11_data_4_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_4_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_4_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_4_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_4_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_4_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_4_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_4_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_4_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_4_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_4_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_4_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_4_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_4_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_4_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_4_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_4_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_4_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_4_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_4_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_4_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_4_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_4_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_4_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_4_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_4_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_4_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_4_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_4_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_4_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_5_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_5_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_5_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_5_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_5_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_5_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_5_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_5_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_5_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_5_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_5_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_5_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_5_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_5_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_5_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_5_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_5_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_5_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_5_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_5_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_5_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_5_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_5_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_5_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_5_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_5_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_5_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_5_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_5_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_5_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_5_cse ) begin
      buffer_bank11_data_5_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_5_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_5_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_5_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_5_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_5_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_5_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_5_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_5_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_5_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_5_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_5_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_5_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_5_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_5_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_5_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_5_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_5_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_5_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_5_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_5_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_5_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_5_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_5_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_5_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_5_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_5_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_5_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_5_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_5_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_6_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_6_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_6_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_6_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_6_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_6_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_6_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_6_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_6_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_6_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_6_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_6_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_6_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_6_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_6_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_6_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_6_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_6_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_6_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_6_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_6_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_6_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_6_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_6_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_6_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_6_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_6_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_6_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_6_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_6_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_6_cse ) begin
      buffer_bank11_data_6_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_6_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_6_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_6_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_6_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_6_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_6_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_6_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_6_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_6_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_6_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_6_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_6_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_6_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_6_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_6_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_6_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_6_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_6_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_6_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_6_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_6_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_6_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_6_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_6_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_6_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_6_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_6_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_6_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_6_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_7_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_7_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_7_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_7_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_7_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_7_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_7_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_7_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_7_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_7_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_7_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_7_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_7_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_7_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_7_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_7_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_7_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_7_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_7_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_7_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_7_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_7_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_7_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_7_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_7_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_7_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_7_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_7_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_7_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_7_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_7_cse ) begin
      buffer_bank11_data_7_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_7_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_7_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_7_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_7_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_7_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_7_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_7_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_7_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_7_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_7_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_7_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_7_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_7_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_7_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_7_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_7_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_7_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_7_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_7_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_7_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_7_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_7_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_7_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_7_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_7_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_7_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_7_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_7_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_7_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_8_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_8_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_8_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_8_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_8_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_8_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_8_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_8_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_8_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_8_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_8_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_8_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_8_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_8_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_8_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_8_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_8_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_8_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_8_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_8_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_8_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_8_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_8_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_8_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_8_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_8_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_8_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_8_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_8_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_8_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_8_cse ) begin
      buffer_bank11_data_8_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_8_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_8_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_8_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_8_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_8_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_8_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_8_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_8_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_8_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_8_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_8_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_8_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_8_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_8_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_8_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_8_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_8_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_8_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_8_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_8_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_8_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_8_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_8_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_8_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_8_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_8_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_8_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_8_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_8_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_9_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_9_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_9_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_9_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_9_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_9_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_9_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_9_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_9_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_9_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_9_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_9_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_9_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_9_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_9_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_9_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_9_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_9_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_9_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_9_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_9_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_9_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_9_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_9_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_9_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_9_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_9_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_9_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_9_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_9_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_9_cse ) begin
      buffer_bank11_data_9_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_9_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_9_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_9_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_9_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_9_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_9_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_9_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_9_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_9_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_9_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_9_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_9_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_9_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_9_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_9_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_9_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_9_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_9_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_9_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_9_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_9_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_9_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_9_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_9_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_9_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_9_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_9_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_9_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_9_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_10_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_10_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_10_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_10_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_10_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_10_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_10_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_10_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_10_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_10_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_10_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_10_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_10_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_10_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_10_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_10_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_10_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_10_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_10_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_10_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_10_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_10_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_10_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_10_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_10_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_10_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_10_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_10_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_10_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_10_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_10_cse ) begin
      buffer_bank11_data_10_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_10_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_10_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_10_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_10_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_10_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_10_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_10_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_10_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_10_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_10_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_10_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_10_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_10_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_10_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_10_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_10_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_10_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_10_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_10_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_10_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_10_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_10_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_10_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_10_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_10_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_10_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_10_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_10_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_10_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_11_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_11_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_11_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_11_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_11_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_11_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_11_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_11_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_11_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_11_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_11_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_11_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_11_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_11_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_11_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_11_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_11_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_11_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_11_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_11_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_11_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_11_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_11_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_11_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_11_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_11_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_11_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_11_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_11_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_11_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_11_cse ) begin
      buffer_bank11_data_11_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_11_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_11_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_11_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_11_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_11_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_11_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_11_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_11_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_11_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_11_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_11_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_11_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_11_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_11_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_11_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_11_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_11_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_11_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_11_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_11_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_11_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_11_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_11_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_11_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_11_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_11_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_11_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_11_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_11_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_12_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_12_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_12_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_12_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_12_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_12_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_12_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_12_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_12_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_12_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_12_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_12_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_12_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_12_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_12_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_12_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_12_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_12_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_12_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_12_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_12_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_12_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_12_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_12_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_12_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_12_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_12_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_12_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_12_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_12_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_12_cse ) begin
      buffer_bank11_data_12_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_12_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_12_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_12_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_12_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_12_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_12_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_12_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_12_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_12_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_12_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_12_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_12_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_12_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_12_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_12_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_12_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_12_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_12_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_12_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_12_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_12_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_12_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_12_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_12_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_12_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_12_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_12_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_12_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_12_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_13_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_13_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_13_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_13_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_13_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_13_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_13_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_13_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_13_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_13_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_13_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_13_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_13_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_13_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_13_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_13_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_13_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_13_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_13_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_13_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_13_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_13_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_13_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_13_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_13_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_13_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_13_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_13_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_13_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_13_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_13_cse ) begin
      buffer_bank11_data_13_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_13_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_13_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_13_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_13_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_13_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_13_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_13_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_13_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_13_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_13_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_13_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_13_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_13_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_13_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_13_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_13_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_13_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_13_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_13_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_13_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_13_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_13_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_13_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_13_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_13_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_13_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_13_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_13_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_13_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_14_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_14_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_14_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_14_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_14_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_14_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_14_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_14_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_14_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_14_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_14_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_14_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_14_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_14_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_14_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_14_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_14_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_14_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_14_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_14_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_14_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_14_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_14_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_14_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_14_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_14_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_14_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_14_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_14_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_14_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_14_cse ) begin
      buffer_bank11_data_14_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_14_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_14_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_14_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_14_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_14_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_14_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_14_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_14_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_14_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_14_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_14_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_14_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_14_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_14_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_14_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_14_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_14_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_14_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_14_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_14_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_14_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_14_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_14_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_14_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_14_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_14_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_14_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_14_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_14_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_15_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_15_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_15_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_15_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_15_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_15_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_15_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_15_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_15_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_15_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_15_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_15_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_15_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_15_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_15_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_15_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_15_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_15_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_15_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_15_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_15_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_15_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_15_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_15_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_15_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_15_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_15_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_15_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_15_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_15_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_15_cse ) begin
      buffer_bank11_data_15_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_15_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_15_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_15_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_15_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_15_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_15_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_15_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_15_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_15_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_15_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_15_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_15_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_15_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_15_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_15_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_15_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_15_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_15_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_15_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_15_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_15_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_15_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_15_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_15_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_15_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_15_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_15_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_15_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_15_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_16_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_16_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_16_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_16_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_16_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_16_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_16_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_16_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_16_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_16_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_16_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_16_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_16_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_16_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_16_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_16_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_16_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_16_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_16_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_16_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_16_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_16_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_16_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_16_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_16_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_16_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_16_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_16_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_16_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_16_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_16_cse ) begin
      buffer_bank11_data_16_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_16_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_16_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_16_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_16_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_16_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_16_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_16_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_16_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_16_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_16_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_16_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_16_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_16_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_16_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_16_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_16_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_16_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_16_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_16_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_16_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_16_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_16_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_16_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_16_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_16_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_16_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_16_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_16_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_16_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_17_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_17_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_17_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_17_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_17_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_17_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_17_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_17_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_17_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_17_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_17_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_17_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_17_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_17_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_17_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_17_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_17_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_17_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_17_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_17_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_17_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_17_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_17_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_17_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_17_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_17_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_17_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_17_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_17_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_17_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_17_cse ) begin
      buffer_bank11_data_17_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_17_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_17_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_17_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_17_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_17_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_17_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_17_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_17_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_17_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_17_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_17_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_17_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_17_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_17_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_17_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_17_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_17_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_17_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_17_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_17_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_17_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_17_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_17_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_17_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_17_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_17_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_17_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_17_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_17_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_18_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_18_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_18_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_18_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_18_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_18_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_18_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_18_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_18_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_18_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_18_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_18_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_18_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_18_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_18_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_18_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_18_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_18_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_18_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_18_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_18_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_18_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_18_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_18_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_18_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_18_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_18_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_18_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_18_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_18_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_18_cse ) begin
      buffer_bank11_data_18_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_18_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_18_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_18_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_18_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_18_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_18_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_18_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_18_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_18_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_18_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_18_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_18_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_18_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_18_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_18_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_18_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_18_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_18_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_18_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_18_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_18_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_18_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_18_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_18_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_18_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_18_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_18_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_18_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_18_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_19_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_19_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_19_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_19_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_19_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_19_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_19_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_19_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_19_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_19_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_19_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_19_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_19_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_19_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_19_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_19_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_19_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_19_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_19_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_19_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_19_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_19_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_19_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_19_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_19_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_19_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_19_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_19_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_19_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_19_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_19_cse ) begin
      buffer_bank11_data_19_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_19_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_19_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_19_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_19_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_19_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_19_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_19_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_19_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_19_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_19_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_19_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_19_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_19_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_19_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_19_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_19_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_19_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_19_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_19_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_19_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_19_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_19_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_19_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_19_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_19_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_19_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_19_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_19_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_19_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_20_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_20_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_20_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_20_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_20_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_20_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_20_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_20_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_20_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_20_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_20_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_20_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_20_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_20_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_20_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_20_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_20_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_20_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_20_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_20_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_20_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_20_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_20_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_20_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_20_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_20_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_20_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_20_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_20_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_20_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_20_cse ) begin
      buffer_bank11_data_20_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_20_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_20_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_20_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_20_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_20_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_20_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_20_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_20_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_20_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_20_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_20_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_20_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_20_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_20_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_20_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_20_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_20_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_20_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_20_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_20_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_20_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_20_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_20_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_20_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_20_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_20_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_20_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_20_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_20_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_21_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_21_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_21_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_21_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_21_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_21_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_21_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_21_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_21_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_21_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_21_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_21_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_21_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_21_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_21_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_21_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_21_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_21_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_21_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_21_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_21_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_21_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_21_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_21_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_21_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_21_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_21_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_21_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_21_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_21_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_21_cse ) begin
      buffer_bank11_data_21_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_21_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_21_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_21_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_21_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_21_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_21_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_21_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_21_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_21_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_21_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_21_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_21_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_21_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_21_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_21_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_21_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_21_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_21_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_21_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_21_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_21_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_21_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_21_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_21_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_21_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_21_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_21_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_21_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_21_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_22_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_22_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_22_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_22_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_22_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_22_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_22_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_22_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_22_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_22_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_22_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_22_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_22_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_22_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_22_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_22_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_22_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_22_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_22_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_22_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_22_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_22_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_22_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_22_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_22_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_22_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_22_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_22_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_22_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_22_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_22_cse ) begin
      buffer_bank11_data_22_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_22_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_22_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_22_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_22_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_22_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_22_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_22_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_22_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_22_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_22_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_22_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_22_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_22_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_22_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_22_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_22_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_22_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_22_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_22_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_22_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_22_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_22_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_22_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_22_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_22_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_22_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_22_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_22_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_22_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_23_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_23_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_23_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_23_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_23_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_23_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_23_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_23_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_23_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_23_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_23_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_23_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_23_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_23_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_23_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_23_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_23_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_23_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_23_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_23_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_23_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_23_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_23_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_23_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_23_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_23_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_23_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_23_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_23_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_23_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_23_cse ) begin
      buffer_bank11_data_23_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_23_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_23_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_23_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_23_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_23_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_23_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_23_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_23_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_23_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_23_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_23_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_23_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_23_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_23_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_23_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_23_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_23_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_23_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_23_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_23_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_23_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_23_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_23_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_23_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_23_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_23_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_23_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_23_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_23_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_24_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_24_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_24_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_24_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_24_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_24_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_24_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_24_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_24_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_24_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_24_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_24_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_24_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_24_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_24_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_24_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_24_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_24_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_24_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_24_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_24_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_24_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_24_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_24_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_24_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_24_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_24_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_24_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_24_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_24_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_24_cse ) begin
      buffer_bank11_data_24_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_24_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_24_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_24_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_24_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_24_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_24_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_24_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_24_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_24_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_24_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_24_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_24_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_24_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_24_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_24_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_24_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_24_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_24_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_24_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_24_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_24_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_24_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_24_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_24_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_24_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_24_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_24_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_24_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_24_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_25_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_25_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_25_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_25_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_25_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_25_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_25_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_25_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_25_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_25_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_25_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_25_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_25_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_25_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_25_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_25_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_25_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_25_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_25_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_25_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_25_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_25_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_25_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_25_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_25_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_25_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_25_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_25_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_25_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_25_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_25_cse ) begin
      buffer_bank11_data_25_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_25_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_25_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_25_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_25_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_25_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_25_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_25_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_25_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_25_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_25_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_25_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_25_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_25_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_25_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_25_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_25_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_25_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_25_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_25_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_25_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_25_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_25_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_25_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_25_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_25_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_25_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_25_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_25_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_25_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_26_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_26_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_26_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_26_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_26_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_26_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_26_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_26_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_26_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_26_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_26_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_26_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_26_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_26_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_26_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_26_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_26_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_26_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_26_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_26_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_26_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_26_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_26_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_26_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_26_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_26_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_26_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_26_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_26_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_26_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_26_cse ) begin
      buffer_bank11_data_26_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_26_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_26_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_26_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_26_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_26_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_26_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_26_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_26_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_26_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_26_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_26_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_26_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_26_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_26_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_26_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_26_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_26_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_26_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_26_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_26_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_26_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_26_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_26_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_26_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_26_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_26_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_26_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_26_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_26_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_27_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_27_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_27_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_27_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_27_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_27_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_27_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_27_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_27_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_27_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_27_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_27_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_27_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_27_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_27_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_27_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_27_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_27_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_27_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_27_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_27_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_27_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_27_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_27_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_27_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_27_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_27_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_27_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_27_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_27_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_27_cse ) begin
      buffer_bank11_data_27_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_27_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_27_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_27_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_27_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_27_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_27_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_27_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_27_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_27_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_27_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_27_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_27_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_27_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_27_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_27_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_27_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_27_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_27_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_27_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_27_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_27_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_27_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_27_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_27_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_27_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_27_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_27_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_27_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_27_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_28_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_28_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_28_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_28_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_28_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_28_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_28_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_28_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_28_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_28_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_28_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_28_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_28_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_28_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_28_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_28_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_28_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_28_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_28_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_28_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_28_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_28_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_28_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_28_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_28_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_28_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_28_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_28_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_28_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_28_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_28_cse ) begin
      buffer_bank11_data_28_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_28_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_28_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_28_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_28_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_28_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_28_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_28_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_28_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_28_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_28_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_28_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_28_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_28_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_28_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_28_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_28_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_28_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_28_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_28_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_28_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_28_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_28_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_28_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_28_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_28_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_28_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_28_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_28_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_28_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_29_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_29_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_29_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_29_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_29_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_29_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_29_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_29_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_29_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_29_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_29_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_29_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_29_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_29_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_29_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_29_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_29_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_29_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_29_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_29_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_29_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_29_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_29_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_29_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_29_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_29_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_29_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_29_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_29_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_29_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_29_cse ) begin
      buffer_bank11_data_29_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_29_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_29_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_29_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_29_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_29_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_29_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_29_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_29_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_29_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_29_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_29_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_29_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_29_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_29_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_29_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_29_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_29_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_29_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_29_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_29_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_29_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_29_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_29_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_29_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_29_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_29_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_29_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_29_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_29_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_30_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_30_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_30_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_30_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_30_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_30_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_30_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_30_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_30_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_30_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_30_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_30_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_30_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_30_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_30_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_30_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_30_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_30_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_30_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_30_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_30_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_30_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_30_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_30_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_30_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_30_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_30_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_30_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_30_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_30_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_30_cse ) begin
      buffer_bank11_data_30_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_30_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_30_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_30_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_30_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_30_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_30_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_30_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_30_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_30_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_30_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_30_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_30_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_30_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_30_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_30_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_30_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_30_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_30_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_30_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_30_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_30_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_30_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_30_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_30_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_30_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_30_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_30_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_30_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_30_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_31_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_31_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_31_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_31_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_31_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_31_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_31_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_31_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_31_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_31_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_31_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_31_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_31_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_31_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_31_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_31_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_31_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_31_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_31_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_31_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_31_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_31_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_31_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_31_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_31_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_31_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_31_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_31_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_31_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_31_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_31_cse ) begin
      buffer_bank11_data_31_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_31_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_31_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_31_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_31_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_31_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_31_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_31_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_31_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_31_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_31_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_31_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_31_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_31_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_31_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_31_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_31_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_31_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_31_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_31_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_31_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_31_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_31_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_31_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_31_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_31_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_31_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_31_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_31_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_31_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_32_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_32_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_32_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_32_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_32_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_32_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_32_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_32_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_32_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_32_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_32_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_32_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_32_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_32_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_32_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_32_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_32_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_32_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_32_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_32_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_32_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_32_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_32_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_32_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_32_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_32_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_32_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_32_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_32_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_32_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_32_cse ) begin
      buffer_bank11_data_32_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_32_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_32_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_32_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_32_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_32_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_32_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_32_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_32_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_32_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_32_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_32_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_32_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_32_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_32_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_32_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_32_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_32_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_32_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_32_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_32_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_32_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_32_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_32_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_32_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_32_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_32_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_32_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_32_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_32_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_33_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_33_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_33_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_33_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_33_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_33_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_33_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_33_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_33_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_33_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_33_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_33_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_33_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_33_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_33_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_33_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_33_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_33_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_33_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_33_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_33_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_33_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_33_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_33_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_33_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_33_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_33_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_33_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_33_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_33_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_33_cse ) begin
      buffer_bank11_data_33_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_33_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_33_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_33_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_33_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_33_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_33_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_33_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_33_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_33_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_33_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_33_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_33_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_33_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_33_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_33_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_33_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_33_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_33_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_33_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_33_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_33_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_33_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_33_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_33_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_33_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_33_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_33_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_33_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_33_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_34_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_34_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_34_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_34_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_34_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_34_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_34_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_34_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_34_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_34_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_34_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_34_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_34_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_34_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_34_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_34_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_34_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_34_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_34_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_34_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_34_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_34_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_34_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_34_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_34_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_34_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_34_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_34_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_34_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_34_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_34_cse ) begin
      buffer_bank11_data_34_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_34_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_34_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_34_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_34_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_34_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_34_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_34_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_34_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_34_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_34_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_34_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_34_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_34_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_34_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_34_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_34_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_34_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_34_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_34_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_34_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_34_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_34_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_34_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_34_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_34_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_34_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_34_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_34_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_34_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_35_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_35_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_35_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_35_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_35_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_35_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_35_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_35_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_35_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_35_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_35_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_35_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_35_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_35_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_35_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_35_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_35_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_35_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_35_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_35_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_35_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_35_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_35_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_35_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_35_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_35_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_35_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_35_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_35_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_35_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_35_cse ) begin
      buffer_bank11_data_35_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_35_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_35_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_35_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_35_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_35_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_35_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_35_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_35_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_35_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_35_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_35_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_35_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_35_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_35_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_35_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_35_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_35_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_35_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_35_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_35_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_35_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_35_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_35_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_35_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_35_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_35_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_35_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_35_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_35_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_36_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_36_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_36_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_36_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_36_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_36_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_36_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_36_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_36_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_36_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_36_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_36_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_36_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_36_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_36_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_36_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_36_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_36_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_36_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_36_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_36_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_36_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_36_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_36_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_36_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_36_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_36_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_36_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_36_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_36_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_36_cse ) begin
      buffer_bank11_data_36_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_36_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_36_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_36_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_36_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_36_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_36_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_36_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_36_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_36_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_36_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_36_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_36_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_36_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_36_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_36_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_36_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_36_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_36_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_36_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_36_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_36_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_36_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_36_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_36_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_36_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_36_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_36_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_36_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_36_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_37_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_37_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_37_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_37_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_37_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_37_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_37_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_37_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_37_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_37_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_37_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_37_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_37_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_37_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_37_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_37_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_37_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_37_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_37_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_37_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_37_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_37_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_37_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_37_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_37_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_37_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_37_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_37_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_37_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_37_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_37_cse ) begin
      buffer_bank11_data_37_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_37_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_37_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_37_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_37_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_37_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_37_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_37_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_37_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_37_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_37_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_37_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_37_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_37_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_37_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_37_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_37_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_37_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_37_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_37_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_37_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_37_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_37_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_37_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_37_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_37_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_37_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_37_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_37_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_37_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_38_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_38_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_38_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_38_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_38_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_38_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_38_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_38_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_38_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_38_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_38_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_38_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_38_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_38_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_38_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_38_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_38_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_38_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_38_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_38_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_38_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_38_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_38_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_38_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_38_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_38_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_38_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_38_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_38_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_38_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_38_cse ) begin
      buffer_bank11_data_38_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_38_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_38_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_38_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_38_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_38_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_38_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_38_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_38_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_38_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_38_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_38_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_38_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_38_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_38_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_38_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_38_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_38_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_38_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_38_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_38_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_38_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_38_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_38_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_38_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_38_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_38_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_38_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_38_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_38_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_39_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_39_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_39_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_39_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_39_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_39_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_39_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_39_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_39_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_39_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_39_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_39_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_39_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_39_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_39_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_39_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_39_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_39_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_39_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_39_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_39_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_39_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_39_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_39_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_39_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_39_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_39_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_39_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_39_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_39_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_39_cse ) begin
      buffer_bank11_data_39_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_39_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_39_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_39_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_39_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_39_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_39_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_39_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_39_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_39_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_39_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_39_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_39_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_39_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_39_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_39_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_39_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_39_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_39_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_39_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_39_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_39_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_39_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_39_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_39_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_39_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_39_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_39_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_39_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_39_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_40_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_40_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_40_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_40_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_40_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_40_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_40_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_40_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_40_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_40_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_40_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_40_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_40_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_40_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_40_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_40_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_40_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_40_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_40_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_40_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_40_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_40_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_40_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_40_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_40_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_40_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_40_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_40_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_40_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_40_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_40_cse ) begin
      buffer_bank11_data_40_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_40_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_40_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_40_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_40_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_40_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_40_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_40_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_40_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_40_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_40_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_40_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_40_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_40_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_40_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_40_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_40_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_40_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_40_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_40_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_40_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_40_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_40_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_40_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_40_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_40_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_40_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_40_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_40_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_40_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_41_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_41_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_41_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_41_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_41_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_41_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_41_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_41_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_41_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_41_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_41_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_41_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_41_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_41_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_41_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_41_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_41_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_41_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_41_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_41_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_41_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_41_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_41_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_41_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_41_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_41_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_41_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_41_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_41_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_41_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_41_cse ) begin
      buffer_bank11_data_41_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_41_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_41_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_41_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_41_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_41_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_41_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_41_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_41_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_41_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_41_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_41_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_41_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_41_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_41_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_41_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_41_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_41_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_41_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_41_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_41_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_41_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_41_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_41_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_41_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_41_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_41_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_41_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_41_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_41_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_42_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_42_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_42_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_42_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_42_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_42_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_42_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_42_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_42_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_42_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_42_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_42_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_42_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_42_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_42_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_42_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_42_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_42_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_42_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_42_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_42_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_42_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_42_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_42_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_42_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_42_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_42_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_42_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_42_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_42_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_42_cse ) begin
      buffer_bank11_data_42_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_42_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_42_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_42_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_42_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_42_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_42_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_42_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_42_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_42_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_42_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_42_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_42_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_42_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_42_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_42_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_42_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_42_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_42_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_42_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_42_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_42_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_42_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_42_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_42_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_42_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_42_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_42_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_42_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_42_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_43_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_43_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_43_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_43_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_43_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_43_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_43_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_43_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_43_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_43_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_43_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_43_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_43_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_43_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_43_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_43_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_43_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_43_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_43_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_43_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_43_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_43_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_43_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_43_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_43_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_43_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_43_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_43_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_43_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_43_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_43_cse ) begin
      buffer_bank11_data_43_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_43_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_43_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_43_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_43_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_43_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_43_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_43_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_43_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_43_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_43_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_43_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_43_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_43_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_43_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_43_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_43_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_43_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_43_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_43_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_43_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_43_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_43_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_43_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_43_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_43_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_43_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_43_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_43_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_43_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_44_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_44_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_44_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_44_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_44_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_44_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_44_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_44_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_44_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_44_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_44_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_44_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_44_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_44_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_44_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_44_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_44_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_44_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_44_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_44_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_44_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_44_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_44_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_44_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_44_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_44_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_44_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_44_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_44_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_44_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_44_cse ) begin
      buffer_bank11_data_44_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_44_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_44_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_44_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_44_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_44_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_44_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_44_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_44_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_44_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_44_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_44_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_44_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_44_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_44_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_44_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_44_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_44_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_44_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_44_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_44_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_44_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_44_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_44_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_44_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_44_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_44_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_44_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_44_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_44_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_45_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_45_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_45_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_45_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_45_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_45_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_45_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_45_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_45_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_45_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_45_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_45_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_45_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_45_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_45_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_45_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_45_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_45_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_45_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_45_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_45_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_45_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_45_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_45_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_45_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_45_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_45_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_45_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_45_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_45_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_45_cse ) begin
      buffer_bank11_data_45_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_45_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_45_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_45_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_45_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_45_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_45_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_45_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_45_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_45_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_45_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_45_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_45_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_45_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_45_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_45_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_45_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_45_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_45_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_45_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_45_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_45_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_45_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_45_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_45_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_45_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_45_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_45_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_45_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_45_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_46_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_46_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_46_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_46_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_46_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_46_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_46_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_46_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_46_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_46_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_46_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_46_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_46_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_46_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_46_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_46_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_46_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_46_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_46_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_46_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_46_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_46_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_46_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_46_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_46_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_46_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_46_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_46_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_46_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_46_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_46_cse ) begin
      buffer_bank11_data_46_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_46_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_46_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_46_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_46_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_46_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_46_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_46_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_46_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_46_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_46_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_46_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_46_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_46_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_46_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_46_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_46_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_46_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_46_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_46_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_46_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_46_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_46_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_46_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_46_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_46_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_46_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_46_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_46_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_46_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_47_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_47_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_47_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_47_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_47_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_47_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_47_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_47_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_47_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_47_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_47_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_47_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_47_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_47_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_47_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_47_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_47_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_47_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_47_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_47_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_47_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_47_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_47_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_47_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_47_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_47_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_47_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_47_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_47_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_47_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_47_cse ) begin
      buffer_bank11_data_47_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_47_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_47_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_47_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_47_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_47_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_47_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_47_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_47_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_47_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_47_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_47_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_47_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_47_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_47_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_47_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_47_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_47_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_47_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_47_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_47_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_47_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_47_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_47_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_47_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_47_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_47_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_47_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_47_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_47_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_48_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_48_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_48_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_48_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_48_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_48_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_48_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_48_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_48_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_48_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_48_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_48_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_48_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_48_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_48_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_48_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_48_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_48_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_48_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_48_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_48_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_48_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_48_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_48_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_48_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_48_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_48_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_48_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_48_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_48_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_48_cse ) begin
      buffer_bank11_data_48_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_48_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_48_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_48_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_48_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_48_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_48_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_48_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_48_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_48_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_48_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_48_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_48_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_48_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_48_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_48_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_48_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_48_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_48_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_48_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_48_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_48_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_48_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_48_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_48_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_48_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_48_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_48_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_48_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_48_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_49_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_49_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_49_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_49_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_49_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_49_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_49_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_49_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_49_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_49_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_49_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_49_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_49_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_49_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_49_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_49_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_49_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_49_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_49_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_49_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_49_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_49_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_49_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_49_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_49_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_49_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_49_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_49_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_49_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_49_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_49_cse ) begin
      buffer_bank11_data_49_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_49_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_49_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_49_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_49_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_49_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_49_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_49_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_49_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_49_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_49_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_49_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_49_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_49_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_49_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_49_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_49_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_49_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_49_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_49_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_49_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_49_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_49_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_49_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_49_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_49_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_49_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_49_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_49_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_49_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_50_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_50_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_50_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_50_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_50_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_50_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_50_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_50_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_50_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_50_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_50_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_50_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_50_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_50_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_50_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_50_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_50_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_50_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_50_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_50_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_50_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_50_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_50_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_50_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_50_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_50_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_50_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_50_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_50_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_50_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_50_cse ) begin
      buffer_bank11_data_50_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_50_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_50_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_50_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_50_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_50_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_50_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_50_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_50_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_50_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_50_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_50_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_50_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_50_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_50_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_50_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_50_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_50_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_50_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_50_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_50_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_50_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_50_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_50_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_50_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_50_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_50_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_50_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_50_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_50_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_51_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_51_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_51_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_51_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_51_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_51_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_51_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_51_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_51_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_51_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_51_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_51_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_51_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_51_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_51_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_51_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_51_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_51_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_51_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_51_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_51_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_51_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_51_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_51_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_51_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_51_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_51_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_51_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_51_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_51_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_51_cse ) begin
      buffer_bank11_data_51_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_51_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_51_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_51_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_51_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_51_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_51_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_51_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_51_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_51_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_51_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_51_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_51_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_51_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_51_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_51_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_51_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_51_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_51_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_51_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_51_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_51_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_51_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_51_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_51_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_51_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_51_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_51_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_51_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_51_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_52_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_52_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_52_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_52_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_52_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_52_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_52_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_52_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_52_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_52_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_52_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_52_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_52_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_52_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_52_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_52_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_52_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_52_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_52_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_52_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_52_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_52_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_52_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_52_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_52_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_52_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_52_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_52_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_52_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_52_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_52_cse ) begin
      buffer_bank11_data_52_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_52_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_52_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_52_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_52_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_52_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_52_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_52_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_52_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_52_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_52_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_52_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_52_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_52_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_52_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_52_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_52_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_52_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_52_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_52_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_52_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_52_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_52_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_52_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_52_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_52_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_52_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_52_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_52_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_52_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_53_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_53_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_53_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_53_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_53_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_53_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_53_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_53_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_53_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_53_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_53_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_53_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_53_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_53_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_53_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_53_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_53_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_53_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_53_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_53_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_53_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_53_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_53_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_53_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_53_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_53_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_53_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_53_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_53_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_53_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_53_cse ) begin
      buffer_bank11_data_53_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_53_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_53_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_53_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_53_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_53_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_53_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_53_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_53_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_53_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_53_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_53_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_53_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_53_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_53_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_53_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_53_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_53_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_53_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_53_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_53_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_53_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_53_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_53_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_53_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_53_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_53_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_53_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_53_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_53_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_54_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_54_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_54_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_54_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_54_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_54_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_54_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_54_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_54_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_54_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_54_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_54_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_54_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_54_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_54_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_54_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_54_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_54_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_54_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_54_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_54_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_54_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_54_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_54_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_54_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_54_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_54_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_54_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_54_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_54_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_54_cse ) begin
      buffer_bank11_data_54_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_54_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_54_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_54_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_54_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_54_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_54_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_54_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_54_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_54_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_54_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_54_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_54_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_54_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_54_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_54_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_54_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_54_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_54_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_54_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_54_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_54_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_54_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_54_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_54_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_54_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_54_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_54_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_54_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_54_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_55_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_55_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_55_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_55_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_55_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_55_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_55_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_55_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_55_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_55_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_55_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_55_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_55_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_55_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_55_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_55_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_55_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_55_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_55_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_55_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_55_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_55_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_55_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_55_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_55_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_55_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_55_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_55_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_55_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_55_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_55_cse ) begin
      buffer_bank11_data_55_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_55_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_55_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_55_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_55_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_55_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_55_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_55_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_55_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_55_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_55_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_55_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_55_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_55_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_55_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_55_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_55_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_55_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_55_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_55_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_55_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_55_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_55_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_55_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_55_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_55_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_55_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_55_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_55_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_55_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_56_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_56_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_56_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_56_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_56_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_56_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_56_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_56_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_56_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_56_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_56_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_56_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_56_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_56_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_56_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_56_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_56_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_56_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_56_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_56_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_56_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_56_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_56_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_56_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_56_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_56_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_56_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_56_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_56_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_56_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_56_cse ) begin
      buffer_bank11_data_56_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_56_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_56_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_56_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_56_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_56_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_56_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_56_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_56_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_56_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_56_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_56_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_56_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_56_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_56_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_56_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_56_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_56_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_56_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_56_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_56_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_56_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_56_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_56_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_56_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_56_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_56_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_56_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_56_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_56_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_57_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_57_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_57_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_57_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_57_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_57_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_57_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_57_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_57_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_57_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_57_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_57_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_57_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_57_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_57_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_57_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_57_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_57_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_57_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_57_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_57_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_57_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_57_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_57_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_57_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_57_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_57_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_57_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_57_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_57_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_57_cse ) begin
      buffer_bank11_data_57_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_57_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_57_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_57_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_57_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_57_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_57_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_57_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_57_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_57_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_57_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_57_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_57_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_57_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_57_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_57_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_57_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_57_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_57_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_57_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_57_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_57_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_57_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_57_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_57_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_57_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_57_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_57_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_57_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_57_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_58_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_58_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_58_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_58_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_58_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_58_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_58_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_58_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_58_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_58_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_58_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_58_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_58_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_58_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_58_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_58_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_58_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_58_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_58_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_58_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_58_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_58_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_58_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_58_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_58_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_58_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_58_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_58_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_58_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_58_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_58_cse ) begin
      buffer_bank11_data_58_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_58_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_58_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_58_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_58_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_58_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_58_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_58_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_58_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_58_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_58_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_58_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_58_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_58_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_58_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_58_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_58_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_58_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_58_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_58_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_58_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_58_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_58_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_58_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_58_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_58_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_58_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_58_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_58_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_58_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_59_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_59_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_59_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_59_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_59_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_59_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_59_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_59_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_59_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_59_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_59_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_59_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_59_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_59_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_59_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_59_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_59_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_59_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_59_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_59_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_59_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_59_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_59_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_59_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_59_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_59_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_59_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_59_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_59_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_59_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_59_cse ) begin
      buffer_bank11_data_59_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_59_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_59_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_59_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_59_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_59_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_59_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_59_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_59_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_59_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_59_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_59_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_59_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_59_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_59_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_59_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_59_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_59_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_59_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_59_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_59_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_59_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_59_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_59_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_59_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_59_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_59_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_59_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_59_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_59_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_60_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_60_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_60_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_60_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_60_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_60_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_60_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_60_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_60_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_60_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_60_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_60_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_60_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_60_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_60_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_60_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_60_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_60_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_60_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_60_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_60_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_60_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_60_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_60_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_60_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_60_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_60_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_60_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_60_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_60_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_60_cse ) begin
      buffer_bank11_data_60_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_60_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_60_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_60_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_60_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_60_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_60_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_60_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_60_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_60_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_60_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_60_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_60_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_60_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_60_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_60_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_60_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_60_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_60_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_60_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_60_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_60_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_60_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_60_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_60_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_60_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_60_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_60_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_60_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_60_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_61_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_61_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_61_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_61_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_61_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_61_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_61_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_61_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_61_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_61_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_61_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_61_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_61_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_61_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_61_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_61_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_61_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_61_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_61_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_61_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_61_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_61_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_61_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_61_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_61_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_61_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_61_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_61_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_61_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_61_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_61_cse ) begin
      buffer_bank11_data_61_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_61_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_61_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_61_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_61_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_61_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_61_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_61_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_61_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_61_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_61_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_61_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_61_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_61_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_61_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_61_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_61_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_61_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_61_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_61_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_61_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_61_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_61_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_61_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_61_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_61_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_61_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_61_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_61_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_61_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank11_data_62_lpi_1 <= 25'b0000000000000000000000000;
      buffer_bank0_data_62_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_62_31_30_lpi_1 <= 2'b00;
      buffer_bank0_data_62_23_12_lpi_1 <= 12'b000000000000;
      buffer_bank10_data_62_29_3_lpi_1 <= 27'b000000000000000000000000000;
      buffer_bank0_data_62_31_24_lpi_1 <= 8'b00000000;
      buffer_bank10_data_62_2_0_lpi_1 <= 3'b000;
      buffer_bank1_data_62_3_0_lpi_1 <= 4'b0000;
      buffer_bank9_data_62_31_8_lpi_1 <= 24'b000000000000000000000000;
      buffer_bank1_data_62_15_4_lpi_1 <= 12'b000000000000;
      buffer_bank9_data_62_7_0_lpi_1 <= 8'b00000000;
      buffer_bank1_data_62_27_16_lpi_1 <= 12'b000000000000;
      buffer_bank8_data_62_31_9_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank1_data_62_31_28_lpi_1 <= 4'b0000;
      buffer_bank8_data_62_8_0_lpi_1 <= 9'b000000000;
      buffer_bank2_data_62_7_0_lpi_1 <= 8'b00000000;
      buffer_bank7_data_62_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_62_19_8_lpi_1 <= 12'b000000000000;
      buffer_bank7_data_62_15_0_lpi_1 <= 16'b0000000000000000;
      buffer_bank2_data_62_31_20_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_62_31_23_lpi_1 <= 9'b000000000;
      buffer_bank3_data_62_11_0_lpi_1 <= 12'b000000000000;
      buffer_bank6_data_62_22_0_lpi_1 <= 23'b00000000000000000000000;
      buffer_bank3_data_62_14_12_lpi_1 <= 3'b000;
      buffer_bank5_data_62_31_30_lpi_1 <= 2'b00;
      buffer_bank5_data_62_29_4_lpi_1 <= 26'b00000000000000000000000000;
      buffer_bank3_data_62_31_16_lpi_1 <= 16'b0000000000000000;
      buffer_bank5_data_62_3_0_lpi_1 <= 4'b0000;
      buffer_bank4_data_62_9_0_lpi_1 <= 10'b0000000000;
      buffer_bank4_data_62_31_10_lpi_1 <= 22'b0000000000000000000000;
    end
    else if ( buffer_bank11_data_and_62_cse ) begin
      buffer_bank11_data_62_lpi_1 <= quads_in_rsci_idat_mxwt[376:352];
      buffer_bank0_data_62_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[11:0];
      buffer_bank10_data_62_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[351:350];
      buffer_bank0_data_62_23_12_lpi_1 <= quads_in_rsci_idat_mxwt[23:12];
      buffer_bank10_data_62_29_3_lpi_1 <= quads_in_rsci_idat_mxwt[349:323];
      buffer_bank0_data_62_31_24_lpi_1 <= quads_in_rsci_idat_mxwt[31:24];
      buffer_bank10_data_62_2_0_lpi_1 <= quads_in_rsci_idat_mxwt[322:320];
      buffer_bank1_data_62_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[35:32];
      buffer_bank9_data_62_31_8_lpi_1 <= quads_in_rsci_idat_mxwt[319:296];
      buffer_bank1_data_62_15_4_lpi_1 <= quads_in_rsci_idat_mxwt[47:36];
      buffer_bank9_data_62_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[295:288];
      buffer_bank1_data_62_27_16_lpi_1 <= quads_in_rsci_idat_mxwt[59:48];
      buffer_bank8_data_62_31_9_lpi_1 <= quads_in_rsci_idat_mxwt[287:265];
      buffer_bank1_data_62_31_28_lpi_1 <= quads_in_rsci_idat_mxwt[63:60];
      buffer_bank8_data_62_8_0_lpi_1 <= quads_in_rsci_idat_mxwt[264:256];
      buffer_bank2_data_62_7_0_lpi_1 <= quads_in_rsci_idat_mxwt[71:64];
      buffer_bank7_data_62_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[255:240];
      buffer_bank2_data_62_19_8_lpi_1 <= quads_in_rsci_idat_mxwt[83:72];
      buffer_bank7_data_62_15_0_lpi_1 <= quads_in_rsci_idat_mxwt[239:224];
      buffer_bank2_data_62_31_20_lpi_1 <= quads_in_rsci_idat_mxwt[95:84];
      buffer_bank6_data_62_31_23_lpi_1 <= quads_in_rsci_idat_mxwt[223:215];
      buffer_bank3_data_62_11_0_lpi_1 <= quads_in_rsci_idat_mxwt[107:96];
      buffer_bank6_data_62_22_0_lpi_1 <= quads_in_rsci_idat_mxwt[214:192];
      buffer_bank3_data_62_14_12_lpi_1 <= quads_in_rsci_idat_mxwt[110:108];
      buffer_bank5_data_62_31_30_lpi_1 <= quads_in_rsci_idat_mxwt[191:190];
      buffer_bank5_data_62_29_4_lpi_1 <= quads_in_rsci_idat_mxwt[189:164];
      buffer_bank3_data_62_31_16_lpi_1 <= quads_in_rsci_idat_mxwt[127:112];
      buffer_bank5_data_62_3_0_lpi_1 <= quads_in_rsci_idat_mxwt[163:160];
      buffer_bank4_data_62_9_0_lpi_1 <= quads_in_rsci_idat_mxwt[137:128];
      buffer_bank4_data_62_31_10_lpi_1 <= quads_in_rsci_idat_mxwt[159:138];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_0_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_9 & for_and_59_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_0_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_1_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_10 & for_and_58_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_1_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_2_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_11 & for_and_57_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_2_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_3_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_12 & for_and_56_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_3_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_4_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_13 & for_and_55_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_4_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_5_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_14 & for_and_54_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_5_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_6_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_15 & for_and_53_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_6_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_7_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_16 & for_and_52_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_7_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_8_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_17 & for_and_51_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_8_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_9_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_18 & for_and_50_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_9_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_10_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_19 & for_and_49_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_10_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_11_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_20 & for_and_48_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_11_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_12_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_21 & for_and_47_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_12_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_13_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_22 & for_and_46_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_13_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_14_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_23 & for_and_45_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_14_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_15_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_24 & for_and_44_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_15_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_16_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_25 & for_and_43_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_16_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_17_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_26 & for_and_41_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_17_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_18_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_27 & for_and_39_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_18_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_19_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_28 & for_and_37_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_19_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_20_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_29 & for_and_35_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_20_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_21_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_30 & for_and_33_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_21_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_22_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_31 & for_and_31_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_22_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_23_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_32 & for_and_29_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_23_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_24_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_33 & for_and_27_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_24_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_25_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_34 & for_and_24_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_25_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_26_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_35 & for_and_21_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_26_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_27_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_36 & for_and_18_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_27_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_28_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_37 & for_and_15_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_28_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_29_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_38 & for_and_11_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_29_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_30_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_39 & for_and_7_tmp & (~ (for_i_6_0_lpi_1_dfm_1_5_0[5]))
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_30_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_31_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_40 & for_and_2_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5:4]==2'b01)
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_31_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_32_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_41 & for_and_59_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_32_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_33_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_42 & for_and_58_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_33_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_34_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_43 & for_and_57_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_34_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_35_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_44 & for_and_56_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_35_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_36_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_45 & for_and_55_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_36_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_37_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_46 & for_and_54_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_37_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_38_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_47 & for_and_53_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_38_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_39_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_48 & for_and_52_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_39_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_40_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_49 & for_and_51_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_40_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_41_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_50 & for_and_50_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_41_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_42_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_51 & for_and_49_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_42_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_43_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_52 & for_and_48_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_43_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_44_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_53 & for_and_47_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_44_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_45_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_54 & for_and_46_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_45_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_46_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_55 & for_and_45_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_46_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_47_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_56 & for_and_44_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_47_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_48_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_57 & for_and_43_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_48_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_49_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_58 & for_and_41_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_49_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_50_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_59 & for_and_39_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_50_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_51_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_60 & for_and_37_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_51_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_52_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_61 & for_and_35_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_52_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_53_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_62 & for_and_33_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_53_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_54_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_63 & for_and_31_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_54_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_55_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_64 & for_and_29_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_55_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_56_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_65 & for_and_27_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_56_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_57_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_66 & for_and_24_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_57_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_58_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_67 & for_and_21_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_58_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_59_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_68 & for_and_18_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_59_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_60_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_69 & for_and_15_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_60_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_61_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_70 & for_and_11_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_61_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      buffer_bank3_data_62_15_lpi_1 <= 1'b0;
    end
    else if ( run_wen & mux_tmp_71 & for_and_7_tmp & (for_i_6_0_lpi_1_dfm_1_5_0[5])
        & (~ or_dcpl_2) ) begin
      buffer_bank3_data_62_15_lpi_1 <= quads_in_rsci_idat_mxwt[111];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_1_for_quad_idx_lpi_1_5_0 <= 6'b000000;
    end
    else if ( run_wen & (~ (mux_10_nl)) & for_1_for_1_and_1_tmp & main_stage_0_2
        ) begin
      for_1_for_quad_idx_lpi_1_5_0 <= operator_7_false_acc_tmp[5:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_1_asn_sft_lpi_1 <= 1'b0;
    end
    else if ( run_wen & (mux_87_nl) & (~(for_1_for_for_1_for_and_1_tmp | or_dcpl_12))
        ) begin
      for_1_asn_sft_lpi_1 <= for_1_for_for_1_for_and_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lfst_exitL_exit_for_1_for_lpi_1 <= 1'b0;
    end
    else if ( run_wen & (~ or_dcpl_12) ) begin
      lfst_exitL_exit_for_1_for_lpi_1 <= ~ for_1_for_1_or_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exitL_exit_for_1_for_lpi_1 <= 1'b0;
    end
    else if ( run_wen & ((~ for_1_for_1_and_2_tmp) | for_1_or_tmp_1) & main_stage_0_2
        ) begin
      exitL_exitL_exit_for_1_for_lpi_1 <= MUX_s_1_2_2((for_for_or_nl), for_1_for_1_or_tmp,
          for_1_for_1_and_1_tmp);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_lpi_1_dfm_56_24 <= 33'b000000000000000000000000000000000;
    end
    else if ( or_1_cse & exitL_exit_for_1_sva & for_1_and_1901_cse ) begin
      paramsIn_crt_lpi_1_dfm_56_24 <= paramsIn_crt_lpi_1_dfm_56_24_mx0;
    end
  end
  assign nl_pixels_in_img_mul_nl = $signed((z_out[11:0])) * $signed(conv_u2s_11_12(paramsIn_crt_lpi_1_dfm_56_24_mx0[10:0]));
  assign pixels_in_img_mul_nl = nl_pixels_in_img_mul_nl[21:0];
  assign for_1_not_3868_nl = ~ mux_89_cse;
  assign nor_100_nl = ~((~ operator_33_true_equal_tmp) | (operator_11_false_2_acc_tmp[11:6]!=6'b000000)
      | (~ mux_tmp_89));
  assign mux_93_nl = MUX_s_1_2_2((nor_100_nl), mux_tmp_89, lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign or_303_nl = exitL_exit_for_1_sva | (~ mux_tmp_93);
  assign nand_12_nl = ~(or_1_cse & mux_tmp_93);
  assign mux_97_nl = MUX_s_1_2_2((or_303_nl), (nand_12_nl), main_stage_0_2);
  assign for_1_for_1_for_not_1_nl = ~ operator_33_true_operator_33_true_or_tmp;
  assign for_for_and_nl = MUX_v_43_2_2(43'b0000000000000000000000000000000000000000000,
      for_1_read_request_lpi_1, (for_1_for_1_for_not_1_nl));
  assign for_1_and_1900_nl = (~ for_1_for_1_if_and_tmp) & for_1_for_if_for_1_for_if_or_tmp
      & (~ for_1_asn_sft_lpi_1_dfm_mx0) & for_1_for_1_and_1_tmp;
  assign nand_11_nl = ~(lfst_exitL_exit_for_1_for_lpi_1 & for_1_asn_sft_lpi_1 & (~
      and_tmp_3));
  assign or_300_nl = operator_43_false_acc_itm_43 | and_tmp_3;
  assign mux_102_nl = MUX_s_1_2_2((nand_11_nl), (or_300_nl), exitL_exitL_exit_for_1_for_lpi_1);
  assign mux_103_nl = MUX_s_1_2_2(or_tmp_183, (mux_102_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign or_299_nl = (~ for_1_for_if_unequal_tmp) | (operator_7_false_acc_tmp[6]);
  assign mux_104_nl = MUX_s_1_2_2(and_tmp_2, (mux_103_nl), or_299_nl);
  assign nand_10_nl = ~(lfst_exitL_exit_for_1_for_lpi_1 & for_1_asn_sft_lpi_1 & (~
      nor_tmp_15));
  assign or_298_nl = operator_43_false_acc_itm_43 | nor_tmp_15;
  assign mux_99_nl = MUX_s_1_2_2((nand_10_nl), (or_298_nl), exitL_exitL_exit_for_1_for_lpi_1);
  assign mux_100_nl = MUX_s_1_2_2((for_acc_1_tmp[6]), (mux_99_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign mux_101_nl = MUX_s_1_2_2(nor_tmp_14, (mux_100_nl), operator_7_false_acc_tmp[6]);
  assign mux_105_nl = MUX_s_1_2_2((mux_104_nl), (mux_101_nl), or_297_cse);
  assign mux_98_nl = MUX_s_1_2_2(and_tmp_2, nor_tmp_14, or_297_cse);
  assign or_292_nl = (~((~ (for_1_read_request_lpi_1[0])) | (~ for_1_if_equal_tmp)
      | (for_1_read_request_lpi_1[7]) | (for_1_read_request_lpi_1[6]) | (for_1_read_request_lpi_1[5])
      | (for_1_read_request_lpi_1[4]) | (for_1_read_request_lpi_1[3]) | (for_1_read_request_lpi_1[36])
      | (for_1_read_request_lpi_1[35]) | (for_1_read_request_lpi_1[34]) | (for_1_read_request_lpi_1[33])
      | (for_1_read_request_lpi_1[2]) | (for_1_read_request_lpi_1[1]) | (for_1_read_request_lpi_1[42])
      | (for_1_read_request_lpi_1[41]) | (for_1_read_request_lpi_1[40]) | (for_1_read_request_lpi_1[39])
      | (for_1_read_request_lpi_1[38]) | (for_1_read_request_lpi_1[37]))) | (lfst_exit_for_1_lpi_1_dfm_1[0]);
  assign mux_106_nl = MUX_s_1_2_2((mux_105_nl), (mux_98_nl), or_292_nl);
  assign or_15_nl = ((operator_33_true_equal_tmp | exitL_exitL_exit_for_1_for_lpi_1
      | (for_acc_1_tmp[6])) & for_1_or_tmp_1) | sfi_exit_for_1_lpi_1 | (~ lfst_exitL_exit_for_1_for_lpi_1)
      | for_1_asn_sft_lpi_1;
  assign or_13_nl = (~ for_1_for_if_unequal_tmp) | (operator_7_false_acc_tmp[6])
      | mux_tmp_2;
  assign mux_8_nl = MUX_s_1_2_2((or_13_nl), or_tmp_5, lfst_exit_for_1_lpi_1_dfm_1[0]);
  assign mux_9_nl = MUX_s_1_2_2((or_15_nl), (mux_8_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign or_11_nl = ((exitL_exitL_exit_for_1_for_lpi_1 | (for_acc_1_tmp[6])) & for_1_or_tmp_1)
      | sfi_exit_for_1_lpi_1 | (~ lfst_exitL_exit_for_1_for_lpi_1) | for_1_asn_sft_lpi_1;
  assign or_9_nl = (operator_7_false_acc_tmp[6]) | mux_tmp_2;
  assign mux_6_nl = MUX_s_1_2_2((or_9_nl), or_tmp_5, lfst_exit_for_1_lpi_1_dfm_1[0]);
  assign mux_7_nl = MUX_s_1_2_2((or_11_nl), (mux_6_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign mux_10_nl = MUX_s_1_2_2((mux_9_nl), (mux_7_nl), or_297_cse);
  assign nor_20_nl = ~(exitL_exitL_exit_for_1_for_lpi_1 | (~ lfst_exitL_exit_for_1_for_lpi_1));
  assign nor_21_nl = ~(exitL_exitL_exit_for_1_for_lpi_1 | (~ lfst_exitL_exit_for_1_for_lpi_1)
      | (for_acc_1_tmp[6]) | and_dcpl_6);
  assign mux_85_nl = MUX_s_1_2_2(lfst_exitL_exit_for_1_for_lpi_1, (nor_21_nl), for_1_or_tmp_1);
  assign nand_8_nl = ~(operator_43_false_acc_itm_43 & or_tmp_161);
  assign mux_82_nl = MUX_s_1_2_2(or_tmp_162, (nand_8_nl), exitL_exitL_exit_for_1_for_lpi_1);
  assign or_164_nl = exitL_exitL_exit_for_1_for_lpi_1 | or_tmp_162;
  assign mux_83_nl = MUX_s_1_2_2((mux_82_nl), (or_164_nl), for_1_or_tmp_1);
  assign nor_22_nl = ~((operator_7_false_acc_tmp[6]) | (mux_83_nl));
  assign nor_23_nl = ~(for_1_or_tmp_1 | exitL_exitL_exit_for_1_for_lpi_1 | (~ lfst_exitL_exit_for_1_for_lpi_1));
  assign mux_84_nl = MUX_s_1_2_2((nor_22_nl), (nor_23_nl), lfst_exit_for_1_lpi_1_dfm_1[0]);
  assign mux_86_nl = MUX_s_1_2_2((mux_85_nl), (mux_84_nl), lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign mux_87_nl = MUX_s_1_2_2((nor_20_nl), (mux_86_nl), main_stage_0_2);
  assign for_for_or_nl = exitL_exitL_exit_for_1_for_lpi_1 | operator_33_true_operator_33_true_or_tmp;
  assign pixels_in_img_mux_2_nl = MUX_v_43_2_2(({32'b11111111111111111111111111111111
      , (paramsIn_crt_lpi_1_dfm_56_24_mx0[32:22])}), for_1_read_request_lpi_1, lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign pixels_in_img_mux_3_nl = MUX_v_11_2_2((~ (paramsIn_crt_lpi_1_dfm_56_24_mx0[21:11])),
      11'b00000000001, lfst_exit_for_1_lpi_1_dfm_1[1]);
  assign nl_acc_nl = ({(pixels_in_img_mux_2_nl) , (~ (lfst_exit_for_1_lpi_1_dfm_1[1]))})
      + conv_u2u_12_44({(pixels_in_img_mux_3_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[43:0];
  assign z_out = readslicef_44_43_1((acc_nl));

  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_64_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [0:0] input_8;
    input [0:0] input_9;
    input [0:0] input_10;
    input [0:0] input_11;
    input [0:0] input_12;
    input [0:0] input_13;
    input [0:0] input_14;
    input [0:0] input_15;
    input [0:0] input_16;
    input [0:0] input_17;
    input [0:0] input_18;
    input [0:0] input_19;
    input [0:0] input_20;
    input [0:0] input_21;
    input [0:0] input_22;
    input [0:0] input_23;
    input [0:0] input_24;
    input [0:0] input_25;
    input [0:0] input_26;
    input [0:0] input_27;
    input [0:0] input_28;
    input [0:0] input_29;
    input [0:0] input_30;
    input [0:0] input_31;
    input [0:0] input_32;
    input [0:0] input_33;
    input [0:0] input_34;
    input [0:0] input_35;
    input [0:0] input_36;
    input [0:0] input_37;
    input [0:0] input_38;
    input [0:0] input_39;
    input [0:0] input_40;
    input [0:0] input_41;
    input [0:0] input_42;
    input [0:0] input_43;
    input [0:0] input_44;
    input [0:0] input_45;
    input [0:0] input_46;
    input [0:0] input_47;
    input [0:0] input_48;
    input [0:0] input_49;
    input [0:0] input_50;
    input [0:0] input_51;
    input [0:0] input_52;
    input [0:0] input_53;
    input [0:0] input_54;
    input [0:0] input_55;
    input [0:0] input_56;
    input [0:0] input_57;
    input [0:0] input_58;
    input [0:0] input_59;
    input [0:0] input_60;
    input [0:0] input_61;
    input [0:0] input_62;
    input [0:0] input_63;
    input [5:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_s_1_64_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_64_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [9:0] input_8;
    input [9:0] input_9;
    input [9:0] input_10;
    input [9:0] input_11;
    input [9:0] input_12;
    input [9:0] input_13;
    input [9:0] input_14;
    input [9:0] input_15;
    input [9:0] input_16;
    input [9:0] input_17;
    input [9:0] input_18;
    input [9:0] input_19;
    input [9:0] input_20;
    input [9:0] input_21;
    input [9:0] input_22;
    input [9:0] input_23;
    input [9:0] input_24;
    input [9:0] input_25;
    input [9:0] input_26;
    input [9:0] input_27;
    input [9:0] input_28;
    input [9:0] input_29;
    input [9:0] input_30;
    input [9:0] input_31;
    input [9:0] input_32;
    input [9:0] input_33;
    input [9:0] input_34;
    input [9:0] input_35;
    input [9:0] input_36;
    input [9:0] input_37;
    input [9:0] input_38;
    input [9:0] input_39;
    input [9:0] input_40;
    input [9:0] input_41;
    input [9:0] input_42;
    input [9:0] input_43;
    input [9:0] input_44;
    input [9:0] input_45;
    input [9:0] input_46;
    input [9:0] input_47;
    input [9:0] input_48;
    input [9:0] input_49;
    input [9:0] input_50;
    input [9:0] input_51;
    input [9:0] input_52;
    input [9:0] input_53;
    input [9:0] input_54;
    input [9:0] input_55;
    input [9:0] input_56;
    input [9:0] input_57;
    input [9:0] input_58;
    input [9:0] input_59;
    input [9:0] input_60;
    input [9:0] input_61;
    input [9:0] input_62;
    input [9:0] input_63;
    input [5:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_10_64_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_64_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [11:0] input_2;
    input [11:0] input_3;
    input [11:0] input_4;
    input [11:0] input_5;
    input [11:0] input_6;
    input [11:0] input_7;
    input [11:0] input_8;
    input [11:0] input_9;
    input [11:0] input_10;
    input [11:0] input_11;
    input [11:0] input_12;
    input [11:0] input_13;
    input [11:0] input_14;
    input [11:0] input_15;
    input [11:0] input_16;
    input [11:0] input_17;
    input [11:0] input_18;
    input [11:0] input_19;
    input [11:0] input_20;
    input [11:0] input_21;
    input [11:0] input_22;
    input [11:0] input_23;
    input [11:0] input_24;
    input [11:0] input_25;
    input [11:0] input_26;
    input [11:0] input_27;
    input [11:0] input_28;
    input [11:0] input_29;
    input [11:0] input_30;
    input [11:0] input_31;
    input [11:0] input_32;
    input [11:0] input_33;
    input [11:0] input_34;
    input [11:0] input_35;
    input [11:0] input_36;
    input [11:0] input_37;
    input [11:0] input_38;
    input [11:0] input_39;
    input [11:0] input_40;
    input [11:0] input_41;
    input [11:0] input_42;
    input [11:0] input_43;
    input [11:0] input_44;
    input [11:0] input_45;
    input [11:0] input_46;
    input [11:0] input_47;
    input [11:0] input_48;
    input [11:0] input_49;
    input [11:0] input_50;
    input [11:0] input_51;
    input [11:0] input_52;
    input [11:0] input_53;
    input [11:0] input_54;
    input [11:0] input_55;
    input [11:0] input_56;
    input [11:0] input_57;
    input [11:0] input_58;
    input [11:0] input_59;
    input [11:0] input_60;
    input [11:0] input_61;
    input [11:0] input_62;
    input [11:0] input_63;
    input [5:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_12_64_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_64_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [5:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_16_64_2 = result;
  end
  endfunction


  function automatic [21:0] MUX_v_22_64_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [21:0] input_2;
    input [21:0] input_3;
    input [21:0] input_4;
    input [21:0] input_5;
    input [21:0] input_6;
    input [21:0] input_7;
    input [21:0] input_8;
    input [21:0] input_9;
    input [21:0] input_10;
    input [21:0] input_11;
    input [21:0] input_12;
    input [21:0] input_13;
    input [21:0] input_14;
    input [21:0] input_15;
    input [21:0] input_16;
    input [21:0] input_17;
    input [21:0] input_18;
    input [21:0] input_19;
    input [21:0] input_20;
    input [21:0] input_21;
    input [21:0] input_22;
    input [21:0] input_23;
    input [21:0] input_24;
    input [21:0] input_25;
    input [21:0] input_26;
    input [21:0] input_27;
    input [21:0] input_28;
    input [21:0] input_29;
    input [21:0] input_30;
    input [21:0] input_31;
    input [21:0] input_32;
    input [21:0] input_33;
    input [21:0] input_34;
    input [21:0] input_35;
    input [21:0] input_36;
    input [21:0] input_37;
    input [21:0] input_38;
    input [21:0] input_39;
    input [21:0] input_40;
    input [21:0] input_41;
    input [21:0] input_42;
    input [21:0] input_43;
    input [21:0] input_44;
    input [21:0] input_45;
    input [21:0] input_46;
    input [21:0] input_47;
    input [21:0] input_48;
    input [21:0] input_49;
    input [21:0] input_50;
    input [21:0] input_51;
    input [21:0] input_52;
    input [21:0] input_53;
    input [21:0] input_54;
    input [21:0] input_55;
    input [21:0] input_56;
    input [21:0] input_57;
    input [21:0] input_58;
    input [21:0] input_59;
    input [21:0] input_60;
    input [21:0] input_61;
    input [21:0] input_62;
    input [21:0] input_63;
    input [5:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_22_64_2 = result;
  end
  endfunction


  function automatic [22:0] MUX_v_23_64_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [22:0] input_2;
    input [22:0] input_3;
    input [22:0] input_4;
    input [22:0] input_5;
    input [22:0] input_6;
    input [22:0] input_7;
    input [22:0] input_8;
    input [22:0] input_9;
    input [22:0] input_10;
    input [22:0] input_11;
    input [22:0] input_12;
    input [22:0] input_13;
    input [22:0] input_14;
    input [22:0] input_15;
    input [22:0] input_16;
    input [22:0] input_17;
    input [22:0] input_18;
    input [22:0] input_19;
    input [22:0] input_20;
    input [22:0] input_21;
    input [22:0] input_22;
    input [22:0] input_23;
    input [22:0] input_24;
    input [22:0] input_25;
    input [22:0] input_26;
    input [22:0] input_27;
    input [22:0] input_28;
    input [22:0] input_29;
    input [22:0] input_30;
    input [22:0] input_31;
    input [22:0] input_32;
    input [22:0] input_33;
    input [22:0] input_34;
    input [22:0] input_35;
    input [22:0] input_36;
    input [22:0] input_37;
    input [22:0] input_38;
    input [22:0] input_39;
    input [22:0] input_40;
    input [22:0] input_41;
    input [22:0] input_42;
    input [22:0] input_43;
    input [22:0] input_44;
    input [22:0] input_45;
    input [22:0] input_46;
    input [22:0] input_47;
    input [22:0] input_48;
    input [22:0] input_49;
    input [22:0] input_50;
    input [22:0] input_51;
    input [22:0] input_52;
    input [22:0] input_53;
    input [22:0] input_54;
    input [22:0] input_55;
    input [22:0] input_56;
    input [22:0] input_57;
    input [22:0] input_58;
    input [22:0] input_59;
    input [22:0] input_60;
    input [22:0] input_61;
    input [22:0] input_62;
    input [22:0] input_63;
    input [5:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_23_64_2 = result;
  end
  endfunction


  function automatic [23:0] MUX_v_24_64_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [23:0] input_2;
    input [23:0] input_3;
    input [23:0] input_4;
    input [23:0] input_5;
    input [23:0] input_6;
    input [23:0] input_7;
    input [23:0] input_8;
    input [23:0] input_9;
    input [23:0] input_10;
    input [23:0] input_11;
    input [23:0] input_12;
    input [23:0] input_13;
    input [23:0] input_14;
    input [23:0] input_15;
    input [23:0] input_16;
    input [23:0] input_17;
    input [23:0] input_18;
    input [23:0] input_19;
    input [23:0] input_20;
    input [23:0] input_21;
    input [23:0] input_22;
    input [23:0] input_23;
    input [23:0] input_24;
    input [23:0] input_25;
    input [23:0] input_26;
    input [23:0] input_27;
    input [23:0] input_28;
    input [23:0] input_29;
    input [23:0] input_30;
    input [23:0] input_31;
    input [23:0] input_32;
    input [23:0] input_33;
    input [23:0] input_34;
    input [23:0] input_35;
    input [23:0] input_36;
    input [23:0] input_37;
    input [23:0] input_38;
    input [23:0] input_39;
    input [23:0] input_40;
    input [23:0] input_41;
    input [23:0] input_42;
    input [23:0] input_43;
    input [23:0] input_44;
    input [23:0] input_45;
    input [23:0] input_46;
    input [23:0] input_47;
    input [23:0] input_48;
    input [23:0] input_49;
    input [23:0] input_50;
    input [23:0] input_51;
    input [23:0] input_52;
    input [23:0] input_53;
    input [23:0] input_54;
    input [23:0] input_55;
    input [23:0] input_56;
    input [23:0] input_57;
    input [23:0] input_58;
    input [23:0] input_59;
    input [23:0] input_60;
    input [23:0] input_61;
    input [23:0] input_62;
    input [23:0] input_63;
    input [5:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_24_64_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_64_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [24:0] input_2;
    input [24:0] input_3;
    input [24:0] input_4;
    input [24:0] input_5;
    input [24:0] input_6;
    input [24:0] input_7;
    input [24:0] input_8;
    input [24:0] input_9;
    input [24:0] input_10;
    input [24:0] input_11;
    input [24:0] input_12;
    input [24:0] input_13;
    input [24:0] input_14;
    input [24:0] input_15;
    input [24:0] input_16;
    input [24:0] input_17;
    input [24:0] input_18;
    input [24:0] input_19;
    input [24:0] input_20;
    input [24:0] input_21;
    input [24:0] input_22;
    input [24:0] input_23;
    input [24:0] input_24;
    input [24:0] input_25;
    input [24:0] input_26;
    input [24:0] input_27;
    input [24:0] input_28;
    input [24:0] input_29;
    input [24:0] input_30;
    input [24:0] input_31;
    input [24:0] input_32;
    input [24:0] input_33;
    input [24:0] input_34;
    input [24:0] input_35;
    input [24:0] input_36;
    input [24:0] input_37;
    input [24:0] input_38;
    input [24:0] input_39;
    input [24:0] input_40;
    input [24:0] input_41;
    input [24:0] input_42;
    input [24:0] input_43;
    input [24:0] input_44;
    input [24:0] input_45;
    input [24:0] input_46;
    input [24:0] input_47;
    input [24:0] input_48;
    input [24:0] input_49;
    input [24:0] input_50;
    input [24:0] input_51;
    input [24:0] input_52;
    input [24:0] input_53;
    input [24:0] input_54;
    input [24:0] input_55;
    input [24:0] input_56;
    input [24:0] input_57;
    input [24:0] input_58;
    input [24:0] input_59;
    input [24:0] input_60;
    input [24:0] input_61;
    input [24:0] input_62;
    input [24:0] input_63;
    input [5:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_25_64_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_64_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input [25:0] input_2;
    input [25:0] input_3;
    input [25:0] input_4;
    input [25:0] input_5;
    input [25:0] input_6;
    input [25:0] input_7;
    input [25:0] input_8;
    input [25:0] input_9;
    input [25:0] input_10;
    input [25:0] input_11;
    input [25:0] input_12;
    input [25:0] input_13;
    input [25:0] input_14;
    input [25:0] input_15;
    input [25:0] input_16;
    input [25:0] input_17;
    input [25:0] input_18;
    input [25:0] input_19;
    input [25:0] input_20;
    input [25:0] input_21;
    input [25:0] input_22;
    input [25:0] input_23;
    input [25:0] input_24;
    input [25:0] input_25;
    input [25:0] input_26;
    input [25:0] input_27;
    input [25:0] input_28;
    input [25:0] input_29;
    input [25:0] input_30;
    input [25:0] input_31;
    input [25:0] input_32;
    input [25:0] input_33;
    input [25:0] input_34;
    input [25:0] input_35;
    input [25:0] input_36;
    input [25:0] input_37;
    input [25:0] input_38;
    input [25:0] input_39;
    input [25:0] input_40;
    input [25:0] input_41;
    input [25:0] input_42;
    input [25:0] input_43;
    input [25:0] input_44;
    input [25:0] input_45;
    input [25:0] input_46;
    input [25:0] input_47;
    input [25:0] input_48;
    input [25:0] input_49;
    input [25:0] input_50;
    input [25:0] input_51;
    input [25:0] input_52;
    input [25:0] input_53;
    input [25:0] input_54;
    input [25:0] input_55;
    input [25:0] input_56;
    input [25:0] input_57;
    input [25:0] input_58;
    input [25:0] input_59;
    input [25:0] input_60;
    input [25:0] input_61;
    input [25:0] input_62;
    input [25:0] input_63;
    input [5:0] sel;
    reg [25:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_26_64_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_64_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input [26:0] input_2;
    input [26:0] input_3;
    input [26:0] input_4;
    input [26:0] input_5;
    input [26:0] input_6;
    input [26:0] input_7;
    input [26:0] input_8;
    input [26:0] input_9;
    input [26:0] input_10;
    input [26:0] input_11;
    input [26:0] input_12;
    input [26:0] input_13;
    input [26:0] input_14;
    input [26:0] input_15;
    input [26:0] input_16;
    input [26:0] input_17;
    input [26:0] input_18;
    input [26:0] input_19;
    input [26:0] input_20;
    input [26:0] input_21;
    input [26:0] input_22;
    input [26:0] input_23;
    input [26:0] input_24;
    input [26:0] input_25;
    input [26:0] input_26;
    input [26:0] input_27;
    input [26:0] input_28;
    input [26:0] input_29;
    input [26:0] input_30;
    input [26:0] input_31;
    input [26:0] input_32;
    input [26:0] input_33;
    input [26:0] input_34;
    input [26:0] input_35;
    input [26:0] input_36;
    input [26:0] input_37;
    input [26:0] input_38;
    input [26:0] input_39;
    input [26:0] input_40;
    input [26:0] input_41;
    input [26:0] input_42;
    input [26:0] input_43;
    input [26:0] input_44;
    input [26:0] input_45;
    input [26:0] input_46;
    input [26:0] input_47;
    input [26:0] input_48;
    input [26:0] input_49;
    input [26:0] input_50;
    input [26:0] input_51;
    input [26:0] input_52;
    input [26:0] input_53;
    input [26:0] input_54;
    input [26:0] input_55;
    input [26:0] input_56;
    input [26:0] input_57;
    input [26:0] input_58;
    input [26:0] input_59;
    input [26:0] input_60;
    input [26:0] input_61;
    input [26:0] input_62;
    input [26:0] input_63;
    input [5:0] sel;
    reg [26:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_27_64_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_64_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [1:0] input_2;
    input [1:0] input_3;
    input [1:0] input_4;
    input [1:0] input_5;
    input [1:0] input_6;
    input [1:0] input_7;
    input [1:0] input_8;
    input [1:0] input_9;
    input [1:0] input_10;
    input [1:0] input_11;
    input [1:0] input_12;
    input [1:0] input_13;
    input [1:0] input_14;
    input [1:0] input_15;
    input [1:0] input_16;
    input [1:0] input_17;
    input [1:0] input_18;
    input [1:0] input_19;
    input [1:0] input_20;
    input [1:0] input_21;
    input [1:0] input_22;
    input [1:0] input_23;
    input [1:0] input_24;
    input [1:0] input_25;
    input [1:0] input_26;
    input [1:0] input_27;
    input [1:0] input_28;
    input [1:0] input_29;
    input [1:0] input_30;
    input [1:0] input_31;
    input [1:0] input_32;
    input [1:0] input_33;
    input [1:0] input_34;
    input [1:0] input_35;
    input [1:0] input_36;
    input [1:0] input_37;
    input [1:0] input_38;
    input [1:0] input_39;
    input [1:0] input_40;
    input [1:0] input_41;
    input [1:0] input_42;
    input [1:0] input_43;
    input [1:0] input_44;
    input [1:0] input_45;
    input [1:0] input_46;
    input [1:0] input_47;
    input [1:0] input_48;
    input [1:0] input_49;
    input [1:0] input_50;
    input [1:0] input_51;
    input [1:0] input_52;
    input [1:0] input_53;
    input [1:0] input_54;
    input [1:0] input_55;
    input [1:0] input_56;
    input [1:0] input_57;
    input [1:0] input_58;
    input [1:0] input_59;
    input [1:0] input_60;
    input [1:0] input_61;
    input [1:0] input_62;
    input [1:0] input_63;
    input [5:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_2_64_2 = result;
  end
  endfunction


  function automatic [32:0] MUX_v_33_2_2;
    input [32:0] input_0;
    input [32:0] input_1;
    input [0:0] sel;
    reg [32:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_33_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_64_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [2:0] input_32;
    input [2:0] input_33;
    input [2:0] input_34;
    input [2:0] input_35;
    input [2:0] input_36;
    input [2:0] input_37;
    input [2:0] input_38;
    input [2:0] input_39;
    input [2:0] input_40;
    input [2:0] input_41;
    input [2:0] input_42;
    input [2:0] input_43;
    input [2:0] input_44;
    input [2:0] input_45;
    input [2:0] input_46;
    input [2:0] input_47;
    input [2:0] input_48;
    input [2:0] input_49;
    input [2:0] input_50;
    input [2:0] input_51;
    input [2:0] input_52;
    input [2:0] input_53;
    input [2:0] input_54;
    input [2:0] input_55;
    input [2:0] input_56;
    input [2:0] input_57;
    input [2:0] input_58;
    input [2:0] input_59;
    input [2:0] input_60;
    input [2:0] input_61;
    input [2:0] input_62;
    input [2:0] input_63;
    input [5:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_3_64_2 = result;
  end
  endfunction


  function automatic [42:0] MUX_v_43_2_2;
    input [42:0] input_0;
    input [42:0] input_1;
    input [0:0] sel;
    reg [42:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_43_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_64_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [3:0] input_2;
    input [3:0] input_3;
    input [3:0] input_4;
    input [3:0] input_5;
    input [3:0] input_6;
    input [3:0] input_7;
    input [3:0] input_8;
    input [3:0] input_9;
    input [3:0] input_10;
    input [3:0] input_11;
    input [3:0] input_12;
    input [3:0] input_13;
    input [3:0] input_14;
    input [3:0] input_15;
    input [3:0] input_16;
    input [3:0] input_17;
    input [3:0] input_18;
    input [3:0] input_19;
    input [3:0] input_20;
    input [3:0] input_21;
    input [3:0] input_22;
    input [3:0] input_23;
    input [3:0] input_24;
    input [3:0] input_25;
    input [3:0] input_26;
    input [3:0] input_27;
    input [3:0] input_28;
    input [3:0] input_29;
    input [3:0] input_30;
    input [3:0] input_31;
    input [3:0] input_32;
    input [3:0] input_33;
    input [3:0] input_34;
    input [3:0] input_35;
    input [3:0] input_36;
    input [3:0] input_37;
    input [3:0] input_38;
    input [3:0] input_39;
    input [3:0] input_40;
    input [3:0] input_41;
    input [3:0] input_42;
    input [3:0] input_43;
    input [3:0] input_44;
    input [3:0] input_45;
    input [3:0] input_46;
    input [3:0] input_47;
    input [3:0] input_48;
    input [3:0] input_49;
    input [3:0] input_50;
    input [3:0] input_51;
    input [3:0] input_52;
    input [3:0] input_53;
    input [3:0] input_54;
    input [3:0] input_55;
    input [3:0] input_56;
    input [3:0] input_57;
    input [3:0] input_58;
    input [3:0] input_59;
    input [3:0] input_60;
    input [3:0] input_61;
    input [3:0] input_62;
    input [3:0] input_63;
    input [5:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_4_64_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_64_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [7:0] input_12;
    input [7:0] input_13;
    input [7:0] input_14;
    input [7:0] input_15;
    input [7:0] input_16;
    input [7:0] input_17;
    input [7:0] input_18;
    input [7:0] input_19;
    input [7:0] input_20;
    input [7:0] input_21;
    input [7:0] input_22;
    input [7:0] input_23;
    input [7:0] input_24;
    input [7:0] input_25;
    input [7:0] input_26;
    input [7:0] input_27;
    input [7:0] input_28;
    input [7:0] input_29;
    input [7:0] input_30;
    input [7:0] input_31;
    input [7:0] input_32;
    input [7:0] input_33;
    input [7:0] input_34;
    input [7:0] input_35;
    input [7:0] input_36;
    input [7:0] input_37;
    input [7:0] input_38;
    input [7:0] input_39;
    input [7:0] input_40;
    input [7:0] input_41;
    input [7:0] input_42;
    input [7:0] input_43;
    input [7:0] input_44;
    input [7:0] input_45;
    input [7:0] input_46;
    input [7:0] input_47;
    input [7:0] input_48;
    input [7:0] input_49;
    input [7:0] input_50;
    input [7:0] input_51;
    input [7:0] input_52;
    input [7:0] input_53;
    input [7:0] input_54;
    input [7:0] input_55;
    input [7:0] input_56;
    input [7:0] input_57;
    input [7:0] input_58;
    input [7:0] input_59;
    input [7:0] input_60;
    input [7:0] input_61;
    input [7:0] input_62;
    input [7:0] input_63;
    input [5:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_8_64_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_64_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [8:0] input_2;
    input [8:0] input_3;
    input [8:0] input_4;
    input [8:0] input_5;
    input [8:0] input_6;
    input [8:0] input_7;
    input [8:0] input_8;
    input [8:0] input_9;
    input [8:0] input_10;
    input [8:0] input_11;
    input [8:0] input_12;
    input [8:0] input_13;
    input [8:0] input_14;
    input [8:0] input_15;
    input [8:0] input_16;
    input [8:0] input_17;
    input [8:0] input_18;
    input [8:0] input_19;
    input [8:0] input_20;
    input [8:0] input_21;
    input [8:0] input_22;
    input [8:0] input_23;
    input [8:0] input_24;
    input [8:0] input_25;
    input [8:0] input_26;
    input [8:0] input_27;
    input [8:0] input_28;
    input [8:0] input_29;
    input [8:0] input_30;
    input [8:0] input_31;
    input [8:0] input_32;
    input [8:0] input_33;
    input [8:0] input_34;
    input [8:0] input_35;
    input [8:0] input_36;
    input [8:0] input_37;
    input [8:0] input_38;
    input [8:0] input_39;
    input [8:0] input_40;
    input [8:0] input_41;
    input [8:0] input_42;
    input [8:0] input_43;
    input [8:0] input_44;
    input [8:0] input_45;
    input [8:0] input_46;
    input [8:0] input_47;
    input [8:0] input_48;
    input [8:0] input_49;
    input [8:0] input_50;
    input [8:0] input_51;
    input [8:0] input_52;
    input [8:0] input_53;
    input [8:0] input_54;
    input [8:0] input_55;
    input [8:0] input_56;
    input [8:0] input_57;
    input [8:0] input_58;
    input [8:0] input_59;
    input [8:0] input_60;
    input [8:0] input_61;
    input [8:0] input_62;
    input [8:0] input_63;
    input [5:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_9_64_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_44_1_43;
    input [43:0] vector;
    reg [43:0] tmp;
  begin
    tmp = vector >> 43;
    readslicef_44_1_43 = tmp[0:0];
  end
  endfunction


  function automatic [42:0] readslicef_44_43_1;
    input [43:0] vector;
    reg [43:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_44_43_1 = tmp[42:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [43:0] conv_u2s_43_44 ;
    input [42:0]  vector ;
  begin
    conv_u2s_43_44 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [43:0] conv_u2u_12_44 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_44 = {{32{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper_run
// ------------------------------------------------------------------


module RenderLooper_run (
  clk, arst_n, render_params_rsc_dat, render_params_rsc_vld, render_params_rsc_rdy,
      render_params_out_rsc_dat, render_params_out_rsc_vld, render_params_out_rsc_rdy,
      loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld, loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [419:0] render_params_rsc_dat;
  input render_params_rsc_vld;
  output render_params_rsc_rdy;
  output [419:0] render_params_out_rsc_dat;
  output render_params_out_rsc_vld;
  input render_params_out_rsc_rdy;
  output [22:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire render_params_rsci_wen_comp;
  wire [419:0] render_params_rsci_idat_mxwt;
  wire render_params_out_rsci_wen_comp;
  reg [419:0] render_params_out_rsci_idat;
  wire loopIndicesOut_rsci_wen_comp;
  reg loopIndicesOut_rsci_idat_22;
  reg [10:0] loopIndicesOut_rsci_idat_21_11;
  wire [11:0] nl_loopIndicesOut_rsci_idat_21_11;
  reg [10:0] loopIndicesOut_rsci_idat_10_0;
  wire [1:0] fsm_output;
  wire for_for_for_for_and_3_tmp;
  wire [11:0] for_acc_1_tmp;
  wire [12:0] nl_for_acc_1_tmp;
  wire operator_11_false_3_equal_tmp;
  wire for_for_for_for_for_for_and_2_tmp;
  wire [11:0] for_for_acc_1_tmp;
  wire [12:0] nl_for_for_acc_1_tmp;
  wire [10:0] for_for_for_acc_1_tmp;
  wire [11:0] nl_for_for_for_acc_1_tmp;
  wire operator_33_true_1_equal_1_tmp;
  wire operator_33_true_1_operator_33_true_1_and_tmp;
  wire [5:0] operator_11_false_2_acc_tmp;
  wire [6:0] nl_operator_11_false_2_acc_tmp;
  wire operator_11_false_equal_tmp;
  wire [9:0] for_for_for_for_and_2_tmp;
  wire for_for_or_tmp;
  wire for_and_1_tmp;
  wire or_tmp;
  wire and_dcpl_2;
  wire or_dcpl_11;
  wire and_dcpl_8;
  reg reg_render_params_rsci_oswt_cse;
  wire loopIndicesOut_and_cse;
  reg reg_loopIndicesOut_rsci_ivld_run_psct_cse;
  wire [10:0] stop_point_height_mux_1_cse;
  wire smp_p_pxl_mux_3_cse;
  wire smp_p_pxl_mux_1_cse;
  reg [9:0] for_for_for_samps_10_0_lpi_1_9_0;
  reg exit_for_lpi_1_dfm_2;
  reg exit_for_for_lpi_1_dfm_3;
  reg exitL_exit_for_sva;
  reg else_unequal_tmp;
  reg [10:0] operator_12_true_return_10_0_lpi_1_dfm;
  reg [10:0] operator_11_false_return_10_0_lpi_1_dfm;
  reg smp_p_pxl_10_lpi_1_dfm_2;
  reg smp_p_pxl_8_lpi_1_dfm_2;
  reg exit_for_for_lpi_1_dfm_1;
  reg exit_for_sva_2;
  reg [10:0] for_fy_11_0_lpi_1_10_0;
  reg [10:0] for_for_fx_11_0_lpi_1_10_0;
  reg smp_p_pxl_6_5_lpi_1_dfm_2_1;
  reg smp_p_pxl_6_5_lpi_1_dfm_2_0;
  wire [10:0] for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0;
  wire else_unequal_tmp_mx0w0;
  wire [10:0] operator_11_false_return_10_0_lpi_1_dfm_mx0;
  wire smp_p_pxl_6_5_lpi_1_dfm_2_1_mx0w0;
  wire smp_p_pxl_6_5_lpi_1_dfm_2_0_mx0w0;
  wire operator_2_false_2_operator_2_false_2_and_mdf_sva_1;
  wire [10:0] for_fy_11_0_lpi_1_dfm_10_0_1;
  wire for_and_ssc_1;
  wire and_42_cse;
  wire nand_7_cse;
  wire or_63_cse;
  wire nor_13_cse;

  wire[10:0] mux_1_nl;
  wire[0:0] and_nl;
  wire[0:0] else_mux_1_nl;
  wire[10:0] operator_12_true_acc_nl;
  wire[11:0] nl_operator_12_true_acc_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] mux_nl;
  wire[0:0] or_50_nl;
  wire[0:0] and_60_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] and_59_nl;
  wire[0:0] for_for_not_13_nl;
  wire[0:0] for_mux_14_nl;
  wire[10:0] operator_11_false_acc_nl;
  wire[11:0] nl_operator_11_false_acc_nl;
  wire[0:0] for_mux_12_nl;
  wire[0:0] for_for_mux_1_nl;
  wire[0:0] for_not_16_nl;
  wire[0:0] for_for_for_for_for_for_for_not_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [22:0] nl_RenderLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat;
  assign nl_RenderLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat =
      {loopIndicesOut_rsci_idat_22 , loopIndicesOut_rsci_idat_21_11 , loopIndicesOut_rsci_idat_10_0};
  RenderLooper_run_render_params_rsci RenderLooper_run_render_params_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsc_dat(render_params_rsc_dat),
      .render_params_rsc_vld(render_params_rsc_vld),
      .render_params_rsc_rdy(render_params_rsc_rdy),
      .run_wen(run_wen),
      .render_params_rsci_oswt(reg_render_params_rsci_oswt_cse),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .render_params_rsci_idat_mxwt(render_params_rsci_idat_mxwt)
    );
  RenderLooper_run_render_params_out_rsci RenderLooper_run_render_params_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_out_rsc_dat(render_params_out_rsc_dat),
      .render_params_out_rsc_vld(render_params_out_rsc_vld),
      .render_params_out_rsc_rdy(render_params_out_rsc_rdy),
      .run_wen(run_wen),
      .render_params_out_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .render_params_out_rsci_wen_comp(render_params_out_rsci_wen_comp),
      .render_params_out_rsci_idat(render_params_out_rsci_idat)
    );
  RenderLooper_run_loopIndicesOut_rsci RenderLooper_run_loopIndicesOut_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesOut_rsci_oswt(reg_loopIndicesOut_rsci_ivld_run_psct_cse),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp),
      .loopIndicesOut_rsci_idat(nl_RenderLooper_run_loopIndicesOut_rsci_inst_loopIndicesOut_rsci_idat[22:0])
    );
  RenderLooper_run_staller RenderLooper_run_staller_inst (
      .run_wen(run_wen),
      .render_params_rsci_wen_comp(render_params_rsci_wen_comp),
      .render_params_out_rsci_wen_comp(render_params_out_rsci_wen_comp),
      .loopIndicesOut_rsci_wen_comp(loopIndicesOut_rsci_wen_comp)
    );
  RenderLooper_run_run_fsm RenderLooper_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign loopIndicesOut_and_cse = run_wen & (~ (fsm_output[0]));
  assign smp_p_pxl_mux_1_cse = MUX_s_1_2_2(smp_p_pxl_8_lpi_1_dfm_2, operator_2_false_2_operator_2_false_2_and_mdf_sva_1,
      exitL_exit_for_sva);
  assign or_63_cse = operator_11_false_equal_tmp | (for_for_acc_1_tmp[11]);
  assign nand_7_cse = ~(or_63_cse & (operator_11_false_3_equal_tmp | (for_acc_1_tmp[11]))
      & (for_for_for_acc_1_tmp[10]));
  assign and_42_cse = nand_7_cse & exitL_exit_for_sva & run_wen;
  assign else_mux_1_nl = MUX_s_1_2_2(else_unequal_tmp_mx0w0, else_unequal_tmp, and_dcpl_8);
  assign and_nl = (~ operator_2_false_2_operator_2_false_2_and_mdf_sva_1) & (else_mux_1_nl)
      & or_tmp;
  assign smp_p_pxl_mux_3_cse = MUX_s_1_2_2(smp_p_pxl_10_lpi_1_dfm_2, (and_nl), exitL_exit_for_sva);
  assign nl_operator_12_true_acc_nl = (~ (render_params_rsci_idat_mxwt[126:116]))
      + (render_params_rsci_idat_mxwt[137:127]);
  assign operator_12_true_acc_nl = nl_operator_12_true_acc_nl[10:0];
  assign stop_point_height_mux_1_cse = MUX_v_11_2_2(operator_12_true_return_10_0_lpi_1_dfm,
      (operator_12_true_acc_nl), exitL_exit_for_sva);
  assign nor_13_cse = ~((for_for_acc_1_tmp[11]) | operator_11_false_equal_tmp);
  assign for_for_not_13_nl = ~ for_for_or_tmp;
  assign for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0 = MUX_v_11_2_2(11'b00000000000, for_for_fx_11_0_lpi_1_10_0,
      (for_for_not_13_nl));
  assign for_mux_14_nl = MUX_s_1_2_2(operator_11_false_3_equal_tmp, exit_for_sva_2,
      or_dcpl_11);
  assign for_for_for_for_and_3_tmp = ((for_acc_1_tmp[11]) | (for_mux_14_nl)) & for_for_for_for_for_for_and_2_tmp;
  assign else_unequal_tmp_mx0w0 = ~((render_params_rsci_idat_mxwt[12:11]==2'b01));
  assign nl_operator_11_false_acc_nl = (render_params_rsci_idat_mxwt[115:105]) +
      11'b11111111111;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[10:0];
  assign operator_11_false_return_10_0_lpi_1_dfm_mx0 = MUX_v_11_2_2(operator_11_false_return_10_0_lpi_1_dfm,
      (operator_11_false_acc_nl), exitL_exit_for_sva);
  assign for_mux_12_nl = MUX_s_1_2_2(smp_p_pxl_6_5_lpi_1_dfm_2_1, (~ else_unequal_tmp_mx0w0),
      for_and_1_tmp);
  assign smp_p_pxl_6_5_lpi_1_dfm_2_1_mx0w0 = (for_mux_12_nl) & (~ for_and_ssc_1);
  assign smp_p_pxl_6_5_lpi_1_dfm_2_0_mx0w0 = (smp_p_pxl_6_5_lpi_1_dfm_2_0 & (~ for_and_1_tmp))
      | for_and_ssc_1;
  assign operator_11_false_3_equal_tmp = (for_fy_11_0_lpi_1_dfm_10_0_1) == (stop_point_height_mux_1_cse);
  assign for_for_mux_1_nl = MUX_s_1_2_2(or_63_cse, exit_for_for_lpi_1_dfm_1, and_dcpl_2);
  assign for_for_for_for_for_for_and_2_tmp = (for_for_mux_1_nl) & ((for_for_for_acc_1_tmp[10])
      | operator_33_true_1_operator_33_true_1_and_tmp);
  assign or_tmp = (render_params_rsci_idat_mxwt[12:11]!=2'b00);
  assign operator_2_false_2_operator_2_false_2_and_mdf_sva_1 = (render_params_rsci_idat_mxwt[12:11]==2'b10);
  assign for_not_16_nl = ~ exitL_exit_for_sva;
  assign for_fy_11_0_lpi_1_dfm_10_0_1 = MUX_v_11_2_2(11'b00000000000, for_fy_11_0_lpi_1_10_0,
      (for_not_16_nl));
  assign operator_33_true_1_operator_33_true_1_and_tmp = (for_for_for_for_and_2_tmp[4:0]==5'b11111)
      & operator_33_true_1_equal_1_tmp & (~ (operator_11_false_2_acc_tmp[5]));
  assign for_for_for_for_for_for_for_not_nl = ~ for_for_or_tmp;
  assign for_for_for_for_and_2_tmp = MUX_v_10_2_2(10'b0000000000, for_for_for_samps_10_0_lpi_1_9_0,
      (for_for_for_for_for_for_for_not_nl));
  assign nl_operator_11_false_2_acc_tmp = ({smp_p_pxl_mux_3_cse , 1'b0 , smp_p_pxl_mux_1_cse
      , 1'b0 , smp_p_pxl_6_5_lpi_1_dfm_2_1_mx0w0 , smp_p_pxl_6_5_lpi_1_dfm_2_0_mx0w0})
      + 6'b111111;
  assign operator_11_false_2_acc_tmp = nl_operator_11_false_2_acc_tmp[5:0];
  assign nl_for_acc_1_tmp = conv_u2s_11_12(for_fy_11_0_lpi_1_dfm_10_0_1) + 12'b000000000001;
  assign for_acc_1_tmp = nl_for_acc_1_tmp[11:0];
  assign nl_for_for_acc_1_tmp = conv_u2s_11_12(for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0)
      + 12'b000000000001;
  assign for_for_acc_1_tmp = nl_for_for_acc_1_tmp[11:0];
  assign operator_11_false_equal_tmp = (for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0) ==
      (operator_11_false_return_10_0_lpi_1_dfm_mx0);
  assign nl_for_for_for_acc_1_tmp = conv_u2s_10_11(for_for_for_for_and_2_tmp) + 11'b00000000001;
  assign for_for_for_acc_1_tmp = nl_for_for_for_acc_1_tmp[10:0];
  assign for_for_or_tmp = exit_for_for_lpi_1_dfm_3 | exit_for_lpi_1_dfm_2 | exitL_exit_for_sva;
  assign for_and_1_tmp = or_tmp & exitL_exit_for_sva;
  assign for_and_ssc_1 = (~ or_tmp) & exitL_exit_for_sva;
  assign operator_33_true_1_equal_1_tmp = (for_for_for_for_and_2_tmp[9:5]) == (operator_11_false_2_acc_tmp[4:0]);
  assign and_dcpl_2 = ~((~(exitL_exit_for_sva | exit_for_for_lpi_1_dfm_3 | exit_for_lpi_1_dfm_2
      | (for_for_for_samps_10_0_lpi_1_9_0[4:0]!=5'b11111) | (operator_11_false_2_acc_tmp[5])
      | (~ operator_33_true_1_equal_1_tmp))) | (for_for_for_acc_1_tmp[10]));
  assign or_dcpl_11 = and_dcpl_2 | nor_13_cse;
  assign and_dcpl_8 = ~((render_params_rsci_idat_mxwt[12:11]!=2'b00));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_render_params_rsci_oswt_cse <= 1'b0;
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_render_params_rsci_oswt_cse <= ~((and_dcpl_2 | nor_13_cse | (~(operator_11_false_3_equal_tmp
          | (for_acc_1_tmp[11])))) & (fsm_output[1]));
      reg_loopIndicesOut_rsci_ivld_run_psct_cse <= fsm_output[1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_10_0 <= 11'b00000000000;
      loopIndicesOut_rsci_idat_22 <= 1'b0;
      exitL_exit_for_sva <= 1'b1;
      smp_p_pxl_6_5_lpi_1_dfm_2_1 <= 1'b0;
      smp_p_pxl_6_5_lpi_1_dfm_2_0 <= 1'b0;
      exit_for_lpi_1_dfm_2 <= 1'b0;
      exit_for_for_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( loopIndicesOut_and_cse ) begin
      loopIndicesOut_rsci_idat_10_0 <= for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0;
      loopIndicesOut_rsci_idat_22 <= operator_33_true_1_operator_33_true_1_and_tmp
          & operator_11_false_3_equal_tmp & operator_11_false_equal_tmp;
      exitL_exit_for_sva <= for_for_for_for_and_3_tmp;
      smp_p_pxl_6_5_lpi_1_dfm_2_1 <= smp_p_pxl_6_5_lpi_1_dfm_2_1_mx0w0;
      smp_p_pxl_6_5_lpi_1_dfm_2_0 <= smp_p_pxl_6_5_lpi_1_dfm_2_0_mx0w0;
      exit_for_lpi_1_dfm_2 <= for_for_for_for_and_3_tmp;
      exit_for_for_lpi_1_dfm_3 <= for_for_for_for_for_for_and_2_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      loopIndicesOut_rsci_idat_21_11 <= 11'b00000000000;
    end
    else if ( run_wen & (~((~(exitL_exit_for_sva | exit_for_for_lpi_1_dfm_3 | exit_for_lpi_1_dfm_2))
        | (fsm_output[0]))) ) begin
      loopIndicesOut_rsci_idat_21_11 <= nl_loopIndicesOut_rsci_idat_21_11[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      render_params_out_rsci_idat <= 420'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~((~ exitL_exit_for_sva) | (fsm_output[0]))) ) begin
      render_params_out_rsci_idat <= render_params_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      else_unequal_tmp <= 1'b0;
    end
    else if ( run_wen & (~(and_dcpl_8 | (~ exitL_exit_for_sva) | (fsm_output[0])))
        ) begin
      else_unequal_tmp <= else_unequal_tmp_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      smp_p_pxl_8_lpi_1_dfm_2 <= 1'b0;
      smp_p_pxl_10_lpi_1_dfm_2 <= 1'b0;
      operator_11_false_return_10_0_lpi_1_dfm <= 11'b00000000000;
      operator_12_true_return_10_0_lpi_1_dfm <= 11'b00000000000;
    end
    else if ( and_42_cse ) begin
      smp_p_pxl_8_lpi_1_dfm_2 <= smp_p_pxl_mux_1_cse;
      smp_p_pxl_10_lpi_1_dfm_2 <= smp_p_pxl_mux_3_cse;
      operator_11_false_return_10_0_lpi_1_dfm <= operator_11_false_return_10_0_lpi_1_dfm_mx0;
      operator_12_true_return_10_0_lpi_1_dfm <= stop_point_height_mux_1_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_for_sva_2 <= 1'b0;
    end
    else if ( run_wen & (~(or_dcpl_11 | (fsm_output[0]))) ) begin
      exit_for_sva_2 <= operator_11_false_3_equal_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_for_for_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( run_wen & (~(and_dcpl_2 | (fsm_output[0]))) ) begin
      exit_for_for_lpi_1_dfm_1 <= or_63_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_for_samps_10_0_lpi_1_9_0 <= 10'b0000000000;
    end
    else if ( run_wen & or_dcpl_11 ) begin
      for_for_for_samps_10_0_lpi_1_9_0 <= MUX_v_10_2_2(({{9{or_63_cse}}, or_63_cse}),
          (for_for_for_acc_1_tmp[9:0]), and_dcpl_2);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_fx_11_0_lpi_1_10_0 <= 11'b00000000000;
    end
    else if ( (mux_2_nl) & run_wen ) begin
      for_for_fx_11_0_lpi_1_10_0 <= MUX_v_11_2_2((for_for_acc_1_tmp[10:0]), for_for_fx_11_0_lpi_1_dfm_10_0_mx0w0,
          and_dcpl_2);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_fy_11_0_lpi_1_10_0 <= 11'b00000000000;
    end
    else if ( (mux_3_nl) & run_wen ) begin
      for_fy_11_0_lpi_1_10_0 <= MUX_v_11_2_2((for_acc_1_tmp[10:0]), for_fy_11_0_lpi_1_dfm_10_0_1,
          or_dcpl_11);
    end
  end
  assign mux_1_nl = MUX_v_11_2_2((render_params_out_rsci_idat[126:116]), (render_params_rsci_idat_mxwt[126:116]),
      exitL_exit_for_sva);
  assign nl_loopIndicesOut_rsci_idat_21_11  = for_fy_11_0_lpi_1_dfm_10_0_1 + (mux_1_nl);
  assign or_50_nl = for_for_or_tmp | (~ or_63_cse);
  assign and_60_nl = (for_for_for_samps_10_0_lpi_1_9_0[4:0]==5'b11111) & (~ (operator_11_false_2_acc_tmp[5]))
      & operator_33_true_1_equal_1_tmp;
  assign mux_nl = MUX_s_1_2_2(for_for_or_tmp, (or_50_nl), and_60_nl);
  assign mux_2_nl = MUX_s_1_2_2((mux_nl), (~ or_63_cse), for_for_for_acc_1_tmp[10]);
  assign and_59_nl = ((~(exit_for_for_lpi_1_dfm_3 | exit_for_lpi_1_dfm_2 | (for_for_for_samps_10_0_lpi_1_9_0[4:0]!=5'b11111)
      | (operator_11_false_2_acc_tmp[5]) | (~ operator_33_true_1_equal_1_tmp))) |
      (for_for_for_acc_1_tmp[10])) & (~(nor_13_cse | (for_acc_1_tmp[11]) | operator_11_false_3_equal_tmp));
  assign mux_3_nl = MUX_s_1_2_2((and_59_nl), nand_7_cse, exitL_exit_for_sva);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration_run
// ------------------------------------------------------------------


module RayGeneration_run (
  clk, arst_n, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld, loopIndicesIn_rsc_rdy,
      paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat, paramsOut_rsc_vld,
      paramsOut_rsc_rdy, rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy, psq_vecMul1_run_mul_cmp_a,
      psq_vecMul1_run_mul_cmp_b, psq_vecMul1_run_mul_cmp_z, psq_vecMul1_run_mul_cmp_1_a,
      psq_vecMul1_run_mul_cmp_1_b, psq_vecMul1_run_mul_cmp_1_z, psq_vecMul1_run_mul_cmp_2_a,
      psq_vecMul1_run_mul_cmp_2_b, psq_vecMul1_run_mul_cmp_2_z, psq_vecMul1_run_mul_cmp_3_a,
      psq_vecMul1_run_mul_cmp_3_b, psq_vecMul1_run_mul_cmp_3_z, psq_vecMul1_run_mul_cmp_4_a,
      psq_vecMul1_run_mul_cmp_4_b, psq_vecMul1_run_mul_cmp_4_z, psq_vecMul1_run_mul_cmp_5_a,
      psq_vecMul1_run_mul_cmp_5_b, psq_vecMul1_run_mul_cmp_5_z
);
  input clk;
  input arst_n;
  input [22:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  input [419:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;
  output [24:0] psq_vecMul1_run_mul_cmp_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_a;
  output [31:0] psq_vecMul1_run_mul_cmp_b;
  input [56:0] psq_vecMul1_run_mul_cmp_z;
  output [24:0] psq_vecMul1_run_mul_cmp_1_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_1_a;
  output [31:0] psq_vecMul1_run_mul_cmp_1_b;
  input [56:0] psq_vecMul1_run_mul_cmp_1_z;
  output [24:0] psq_vecMul1_run_mul_cmp_2_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_2_a;
  output [31:0] psq_vecMul1_run_mul_cmp_2_b;
  input [56:0] psq_vecMul1_run_mul_cmp_2_z;
  output [24:0] psq_vecMul1_run_mul_cmp_3_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_3_a;
  output [31:0] psq_vecMul1_run_mul_cmp_3_b;
  input [56:0] psq_vecMul1_run_mul_cmp_3_z;
  output [24:0] psq_vecMul1_run_mul_cmp_4_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_4_a;
  output [31:0] psq_vecMul1_run_mul_cmp_4_b;
  input [56:0] psq_vecMul1_run_mul_cmp_4_z;
  output [24:0] psq_vecMul1_run_mul_cmp_5_a;
  reg [24:0] psq_vecMul1_run_mul_cmp_5_a;
  output [31:0] psq_vecMul1_run_mul_cmp_5_b;
  input [56:0] psq_vecMul1_run_mul_cmp_5_z;


  // Interconnect Declarations
  wire run_wen;
  wire loopIndicesIn_rsci_wen_comp;
  wire [22:0] loopIndicesIn_rsci_idat_mxwt;
  wire paramsIn_rsci_wen_comp;
  wire [373:0] paramsIn_rsci_idat_mxwt;
  wire paramsOut_rsci_wen_comp;
  wire rayOut_rsci_wen_comp;
  wire [24:0] psq_vecMul1_run_mul_cmp_z_oreg;
  wire [24:0] psq_vecMul1_run_mul_cmp_1_z_oreg;
  wire [24:0] psq_vecMul1_run_mul_cmp_2_z_oreg;
  wire [24:0] psq_vecMul1_run_mul_cmp_3_z_oreg;
  wire [24:0] psq_vecMul1_run_mul_cmp_4_z_oreg;
  wire [24:0] psq_vecMul1_run_mul_cmp_5_z_oreg;
  reg paramsOut_rsci_idat_92;
  reg [80:0] paramsOut_rsci_idat_91_11;
  reg [10:0] paramsOut_rsci_idat_10_0;
  reg [10:0] rayOut_rsci_idat_164_154;
  wire [11:0] nl_rayOut_rsci_idat_164_154;
  reg [21:0] rayOut_rsci_idat_153_132;
  reg [10:0] rayOut_rsci_idat_130_120;
  wire [11:0] nl_rayOut_rsci_idat_130_120;
  reg [21:0] rayOut_rsci_idat_119_98;
  reg [10:0] rayOut_rsci_idat_96_86;
  wire [11:0] nl_rayOut_rsci_idat_96_86;
  reg [21:0] rayOut_rsci_idat_85_64;
  reg [10:0] rayOut_rsci_idat_62_52;
  reg [10:0] rayOut_rsci_idat_41_31;
  reg [10:0] rayOut_rsci_idat_20_10;
  reg psq_run_py_not_2;
  reg psq_rand_val2_run_x3_30_sva;
  reg psq_rand_val2_run_x3_29_sva;
  reg psq_rand_val2_run_x3_28_sva;
  reg psq_rand_val2_run_x3_27_sva;
  reg psq_rand_val2_run_x3_26_sva;
  reg psq_rand_val2_run_x3_25_sva;
  reg psq_rand_val2_run_x3_24_sva;
  reg psq_rand_val2_run_x3_23_sva;
  reg psq_rand_val2_run_x3_22_sva;
  reg psq_rand_val2_run_x3_21_sva;
  reg psq_rand_val2_run_x3_20_sva;
  reg psq_rand_val2_run_x3_19_sva;
  reg psq_rand_val2_run_x3_18_sva;
  reg psq_rand_val2_run_x3_17_sva;
  reg psq_rand_val2_run_x3_16_sva;
  reg psq_rand_val2_run_x3_15_sva;
  reg psq_rand_val2_run_x3_14_sva;
  reg psq_rand_val2_run_x3_13_sva;
  reg psq_rand_val2_run_x3_12_sva;
  reg psq_rand_val2_run_x3_11_sva;
  reg psq_rand_val2_run_x3_10_sva;
  reg psq_rand_val2_run_x3_9_sva;
  reg psq_rand_val2_run_x3_8_sva;
  reg psq_rand_val2_run_x3_7_sva;
  reg psq_rand_val2_run_x3_6_sva;
  reg psq_rand_val2_run_x3_5_sva;
  reg psq_rand_val2_run_x2_4_sva;
  reg psq_rand_val2_run_x2_3_sva;
  reg psq_rand_val2_run_x2_2_sva;
  reg psq_rand_val2_run_x2_1_sva;
  reg psq_rand_val2_run_x2_0_sva;
  reg psq_run_px_not_3;
  reg psq_rand_val_run_x3_30_sva;
  reg psq_rand_val_run_x3_29_sva;
  reg psq_rand_val_run_x3_28_sva;
  reg psq_rand_val_run_x3_27_sva;
  reg psq_rand_val_run_x3_26_sva;
  reg psq_rand_val_run_x3_25_sva;
  reg psq_rand_val_run_x3_24_sva;
  reg psq_rand_val_run_x3_23_sva;
  reg psq_rand_val_run_x3_22_sva;
  reg psq_rand_val_run_x3_21_sva;
  reg psq_rand_val_run_x3_20_sva;
  reg psq_rand_val_run_x3_19_sva;
  reg psq_rand_val_run_x3_18_sva;
  reg psq_rand_val_run_x3_17_sva;
  reg psq_rand_val_run_x3_16_sva;
  reg psq_rand_val_run_x3_15_sva;
  reg psq_rand_val_run_x3_14_sva;
  reg psq_rand_val_run_x3_13_sva;
  reg psq_rand_val_run_x3_12_sva;
  reg psq_rand_val_run_x3_11_sva;
  reg psq_rand_val_run_x3_10_sva;
  reg psq_rand_val_run_x3_9_sva;
  reg psq_rand_val_run_x3_8_sva;
  reg psq_rand_val_run_x3_7_sva;
  reg psq_rand_val_run_x3_6_sva;
  reg psq_rand_val_run_x3_5_sva;
  reg psq_rand_val_run_x2_4_sva;
  reg psq_rand_val_run_x2_3_sva;
  reg psq_rand_val_run_x2_2_sva;
  reg psq_rand_val_run_x2_1_sva;
  reg psq_rand_val_run_x2_0_sva;
  wire [1:0] fsm_output;
  wire rayOut_and_cse;
  reg reg_rayOut_rsci_ivld_run_psct_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire state2_and_cse;
  reg main_stage_0_4;
  wire and_itm;
  wire and_132_itm;
  reg state1_15_sva;
  reg state1_16_sva;
  reg state1_14_sva;
  reg state1_17_sva;
  reg state1_13_sva;
  reg state1_18_sva;
  reg state1_12_sva;
  reg state1_19_sva;
  reg state1_11_sva;
  reg state1_20_sva;
  reg state1_10_sva;
  reg state1_21_sva;
  reg state1_9_sva;
  reg state1_22_sva;
  reg state1_8_sva;
  reg state1_23_sva;
  reg state1_7_sva;
  reg state1_24_sva;
  reg state1_6_sva;
  reg state1_25_sva;
  reg state1_5_sva;
  reg state1_26_sva;
  reg state1_4_sva;
  reg state1_27_sva;
  reg state1_3_sva;
  reg state1_28_sva;
  reg state1_2_sva;
  reg state1_29_sva;
  reg state1_1_sva;
  reg state1_30_sva;
  reg state1_0_sva;
  reg state1_31_sva;
  reg state2_15_sva;
  reg state2_16_sva;
  reg state2_14_sva;
  reg state2_17_sva;
  reg state2_13_sva;
  reg state2_18_sva;
  reg state2_12_sva;
  reg state2_19_sva;
  reg state2_11_sva;
  reg state2_20_sva;
  reg state2_10_sva;
  reg state2_21_sva;
  reg state2_9_sva;
  reg state2_22_sva;
  reg state2_8_sva;
  reg state2_23_sva;
  reg state2_7_sva;
  reg state2_24_sva;
  reg state2_6_sva;
  reg state2_25_sva;
  reg state2_5_sva;
  reg state2_26_sva;
  reg state2_4_sva;
  reg state2_27_sva;
  reg state2_3_sva;
  reg state2_28_sva;
  reg state2_2_sva;
  reg state2_29_sva;
  reg state2_1_sva;
  reg state2_30_sva;
  reg state2_0_sva;
  reg state2_31_sva;
  reg main_stage_0_2;
  reg main_stage_0_3;
  reg [32:0] deltUMul_run_mul_itm_1;
  wire signed [36:0] nl_deltUMul_run_mul_itm_1;
  reg [32:0] deltVMul_run_mul_itm_1;
  wire signed [36:0] nl_deltVMul_run_mul_itm_1;
  reg [32:0] deltAdd_run_acc_5_itm_1;
  wire [33:0] nl_deltAdd_run_acc_5_itm_1;
  reg [32:0] deltAdd_run_acc_5_itm_2;
  reg [32:0] deltAdd_run_acc_itm_1;
  wire [33:0] nl_deltAdd_run_acc_itm_1;
  reg [32:0] deltUMul_run_mul_1_itm_1;
  wire signed [36:0] nl_deltUMul_run_mul_1_itm_1;
  reg [32:0] deltVMul_run_mul_1_itm_1;
  wire signed [36:0] nl_deltVMul_run_mul_1_itm_1;
  reg [32:0] deltAdd_run_acc_7_itm_1;
  wire [33:0] nl_deltAdd_run_acc_7_itm_1;
  reg [32:0] deltAdd_run_acc_7_itm_2;
  reg [32:0] deltAdd_run_acc_6_itm_1;
  wire [33:0] nl_deltAdd_run_acc_6_itm_1;
  reg [32:0] deltUMul_run_mul_2_itm_1;
  wire signed [36:0] nl_deltUMul_run_mul_2_itm_1;
  reg [32:0] deltVMul_run_mul_2_itm_1;
  wire signed [36:0] nl_deltVMul_run_mul_2_itm_1;
  reg [32:0] deltAdd_run_acc_9_itm_1;
  wire [33:0] nl_deltAdd_run_acc_9_itm_1;
  reg [32:0] deltAdd_run_acc_9_itm_2;
  reg [32:0] deltAdd_run_acc_8_itm_1;
  wire [33:0] nl_deltAdd_run_acc_8_itm_1;
  reg loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_1;
  reg loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_2;
  reg loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_3;
  reg [131:0] paramsIn_crt_sva_1_269_138;
  reg [80:0] paramsIn_crt_sva_1_93_13;
  reg [10:0] paramsIn_crt_sva_1_10_0;
  reg [131:0] paramsIn_crt_sva_2_269_138;
  reg [80:0] paramsIn_crt_sva_2_93_13;
  reg [10:0] paramsIn_crt_sva_2_10_0;
  reg [32:0] paramsIn_crt_sva_3_170_138;
  reg [80:0] paramsIn_crt_sva_3_93_13;
  reg [10:0] paramsIn_crt_sva_3_10_0;
  wire psq_rand_val2_run_x2_0_sva_4;
  wire psq_rand_val2_run_x2_1_sva_4;
  wire psq_rand_val2_run_x2_2_sva_4;
  wire psq_rand_val2_run_x2_3_sva_4;
  wire psq_rand_val2_run_x2_4_sva_4;
  wire psq_rand_val2_run_x3_5_sva_4;
  wire psq_rand_val2_run_x3_6_sva_4;
  wire psq_rand_val2_run_x3_7_sva_4;
  wire psq_rand_val2_run_x3_8_sva_4;
  wire psq_rand_val2_run_x3_9_sva_4;
  wire psq_rand_val2_run_x3_10_sva_4;
  wire psq_rand_val2_run_x3_11_sva_4;
  wire psq_rand_val2_run_x3_12_sva_4;
  wire psq_rand_val2_run_x3_13_sva_4;
  wire psq_rand_val2_run_x3_14_sva_4;
  wire psq_rand_val2_run_x3_15_sva_4;
  wire psq_rand_val2_run_x3_16_sva_4;
  wire psq_rand_val2_run_x3_17_sva_4;
  wire psq_rand_val2_run_x3_18_sva_4;
  wire psq_rand_val2_run_x3_19_sva_4;
  wire psq_rand_val2_run_x3_20_sva_4;
  wire psq_rand_val2_run_x3_21_sva_4;
  wire psq_rand_val2_run_x3_22_sva_4;
  wire psq_rand_val2_run_x3_23_sva_4;
  wire psq_rand_val2_run_x3_24_sva_4;
  wire psq_rand_val2_run_x3_25_sva_4;
  wire psq_rand_val2_run_x3_26_sva_4;
  wire psq_rand_val2_run_x3_27_sva_4;
  wire psq_rand_val2_run_x3_28_sva_4;
  wire psq_rand_val2_run_x3_29_sva_4;
  wire psq_rand_val2_run_x3_30_sva_4;
  wire psq_rand_val_run_x2_0_sva_4;
  wire psq_rand_val_run_x2_1_sva_4;
  wire psq_rand_val_run_x2_2_sva_4;
  wire psq_rand_val_run_x2_3_sva_4;
  wire psq_rand_val_run_x2_4_sva_4;
  wire psq_rand_val_run_x3_5_sva_4;
  wire psq_rand_val_run_x3_6_sva_4;
  wire psq_rand_val_run_x3_7_sva_4;
  wire psq_rand_val_run_x3_8_sva_4;
  wire psq_rand_val_run_x3_9_sva_4;
  wire psq_rand_val_run_x3_10_sva_4;
  wire psq_rand_val_run_x3_11_sva_4;
  wire psq_rand_val_run_x3_12_sva_4;
  wire psq_rand_val_run_x3_13_sva_4;
  wire psq_rand_val_run_x3_14_sva_4;
  wire psq_rand_val_run_x3_15_sva_4;
  wire psq_rand_val_run_x3_16_sva_4;
  wire psq_rand_val_run_x3_17_sva_4;
  wire psq_rand_val_run_x3_18_sva_4;
  wire psq_rand_val_run_x3_19_sva_4;
  wire psq_rand_val_run_x3_20_sva_4;
  wire psq_rand_val_run_x3_21_sva_4;
  wire psq_rand_val_run_x3_22_sva_4;
  wire psq_rand_val_run_x3_23_sva_4;
  wire psq_rand_val_run_x3_24_sva_4;
  wire psq_rand_val_run_x3_25_sva_4;
  wire psq_rand_val_run_x3_26_sva_4;
  wire psq_rand_val_run_x3_27_sva_4;
  wire psq_rand_val_run_x3_28_sva_4;
  wire psq_rand_val_run_x3_29_sva_4;
  wire psq_rand_val_run_x3_30_sva_4;
  wire [32:0] sampleAdd_run_acc_4_psp_sva_1;
  wire [33:0] nl_sampleAdd_run_acc_4_psp_sva_1;
  wire [32:0] sampleAdd_run_acc_3_psp_sva_1;
  wire [33:0] nl_sampleAdd_run_acc_3_psp_sva_1;
  wire [32:0] sampleAdd_run_acc_psp_sva_1;
  wire [33:0] nl_sampleAdd_run_acc_psp_sva_1;
  wire xor_cse;
  wire xor_cse_1;
  wire xor_cse_2;
  wire xor_cse_3;
  wire xor_cse_4;
  wire xor_cse_5;
  wire xor_cse_6;
  wire xor_cse_7;
  wire xor_cse_8;
  wire xor_cse_10;
  wire xor_cse_11;
  wire xor_cse_12;
  wire xor_cse_13;
  wire xor_cse_14;
  wire xor_cse_15;
  wire xor_cse_16;
  wire xor_cse_17;
  wire xor_cse_18;
  wire xor_cse_20;
  wire xor_cse_21;

  wire[24:0] psq_run_acc_2_nl;
  wire[25:0] nl_psq_run_acc_2_nl;
  wire[24:0] psq_run_acc_1_nl;
  wire[25:0] nl_psq_run_acc_1_nl;
  wire[24:0] psq_run_acc_nl;
  wire[25:0] nl_psq_run_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [92:0] nl_RayGeneration_run_paramsOut_rsci_inst_paramsOut_rsci_idat;
  assign nl_RayGeneration_run_paramsOut_rsci_inst_paramsOut_rsci_idat = {paramsOut_rsci_idat_92
      , paramsOut_rsci_idat_91_11 , paramsOut_rsci_idat_10_0};
  wire [165:0] nl_RayGeneration_run_rayOut_rsci_inst_rayOut_rsci_idat;
  assign nl_RayGeneration_run_rayOut_rsci_inst_rayOut_rsci_idat = {1'b1 , rayOut_rsci_idat_164_154
      , rayOut_rsci_idat_153_132 , 1'b0 , rayOut_rsci_idat_130_120 , rayOut_rsci_idat_119_98
      , 1'b0 , rayOut_rsci_idat_96_86 , rayOut_rsci_idat_85_64 , 1'b0 , rayOut_rsci_idat_62_52
      , 10'b0000000000 , rayOut_rsci_idat_41_31 , 10'b0000000000 , rayOut_rsci_idat_20_10
      , 10'b0000000000};
  RayGeneration_run_loopIndicesIn_rsci RayGeneration_run_loopIndicesIn_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .run_wen(run_wen),
      .loopIndicesIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .loopIndicesIn_rsci_idat_mxwt(loopIndicesIn_rsci_idat_mxwt)
    );
  RayGeneration_run_paramsIn_rsci RayGeneration_run_paramsIn_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  RayGeneration_run_paramsOut_rsci RayGeneration_run_paramsOut_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(reg_rayOut_rsci_ivld_run_psct_cse),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_idat(nl_RayGeneration_run_paramsOut_rsci_inst_paramsOut_rsci_idat[92:0])
    );
  RayGeneration_run_rayOut_rsci RayGeneration_run_rayOut_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rayOut_rsc_dat(rayOut_rsc_dat),
      .rayOut_rsc_vld(rayOut_rsc_vld),
      .rayOut_rsc_rdy(rayOut_rsc_rdy),
      .run_wen(run_wen),
      .rayOut_rsci_oswt(reg_rayOut_rsci_ivld_run_psct_cse),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp),
      .rayOut_rsci_idat(nl_RayGeneration_run_rayOut_rsci_inst_rayOut_rsci_idat[165:0])
    );
  RayGeneration_run_wait_dp RayGeneration_run_wait_dp_inst (
      .clk(clk),
      .arst_n(arst_n),
      .psq_vecMul1_run_mul_cmp_z(psq_vecMul1_run_mul_cmp_z),
      .psq_vecMul1_run_mul_cmp_1_z(psq_vecMul1_run_mul_cmp_1_z),
      .psq_vecMul1_run_mul_cmp_2_z(psq_vecMul1_run_mul_cmp_2_z),
      .psq_vecMul1_run_mul_cmp_3_z(psq_vecMul1_run_mul_cmp_3_z),
      .psq_vecMul1_run_mul_cmp_4_z(psq_vecMul1_run_mul_cmp_4_z),
      .psq_vecMul1_run_mul_cmp_5_z(psq_vecMul1_run_mul_cmp_5_z),
      .run_wen(run_wen),
      .psq_vecMul1_run_mul_cmp_z_oreg(psq_vecMul1_run_mul_cmp_z_oreg),
      .psq_vecMul1_run_mul_cmp_1_z_oreg(psq_vecMul1_run_mul_cmp_1_z_oreg),
      .psq_vecMul1_run_mul_cmp_2_z_oreg(psq_vecMul1_run_mul_cmp_2_z_oreg),
      .psq_vecMul1_run_mul_cmp_3_z_oreg(psq_vecMul1_run_mul_cmp_3_z_oreg),
      .psq_vecMul1_run_mul_cmp_4_z_oreg(psq_vecMul1_run_mul_cmp_4_z_oreg),
      .psq_vecMul1_run_mul_cmp_5_z_oreg(psq_vecMul1_run_mul_cmp_5_z_oreg)
    );
  RayGeneration_run_staller RayGeneration_run_staller_inst (
      .run_wen(run_wen),
      .loopIndicesIn_rsci_wen_comp(loopIndicesIn_rsci_wen_comp),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp)
    );
  RayGeneration_run_run_fsm RayGeneration_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign psq_vecMul1_run_mul_cmp_5_b = {psq_run_py_not_2 , psq_rand_val2_run_x3_30_sva
      , psq_rand_val2_run_x3_29_sva , psq_rand_val2_run_x3_28_sva , psq_rand_val2_run_x3_27_sva
      , psq_rand_val2_run_x3_26_sva , psq_rand_val2_run_x3_25_sva , psq_rand_val2_run_x3_24_sva
      , psq_rand_val2_run_x3_23_sva , psq_rand_val2_run_x3_22_sva , psq_rand_val2_run_x3_21_sva
      , psq_rand_val2_run_x3_20_sva , psq_rand_val2_run_x3_19_sva , psq_rand_val2_run_x3_18_sva
      , psq_rand_val2_run_x3_17_sva , psq_rand_val2_run_x3_16_sva , psq_rand_val2_run_x3_15_sva
      , psq_rand_val2_run_x3_14_sva , psq_rand_val2_run_x3_13_sva , psq_rand_val2_run_x3_12_sva
      , psq_rand_val2_run_x3_11_sva , psq_rand_val2_run_x3_10_sva , psq_rand_val2_run_x3_9_sva
      , psq_rand_val2_run_x3_8_sva , psq_rand_val2_run_x3_7_sva , psq_rand_val2_run_x3_6_sva
      , psq_rand_val2_run_x3_5_sva , psq_rand_val2_run_x2_4_sva , psq_rand_val2_run_x2_3_sva
      , psq_rand_val2_run_x2_2_sva , psq_rand_val2_run_x2_1_sva , psq_rand_val2_run_x2_0_sva};
  assign psq_vecMul1_run_mul_cmp_4_b = {psq_run_px_not_3 , psq_rand_val_run_x3_30_sva
      , psq_rand_val_run_x3_29_sva , psq_rand_val_run_x3_28_sva , psq_rand_val_run_x3_27_sva
      , psq_rand_val_run_x3_26_sva , psq_rand_val_run_x3_25_sva , psq_rand_val_run_x3_24_sva
      , psq_rand_val_run_x3_23_sva , psq_rand_val_run_x3_22_sva , psq_rand_val_run_x3_21_sva
      , psq_rand_val_run_x3_20_sva , psq_rand_val_run_x3_19_sva , psq_rand_val_run_x3_18_sva
      , psq_rand_val_run_x3_17_sva , psq_rand_val_run_x3_16_sva , psq_rand_val_run_x3_15_sva
      , psq_rand_val_run_x3_14_sva , psq_rand_val_run_x3_13_sva , psq_rand_val_run_x3_12_sva
      , psq_rand_val_run_x3_11_sva , psq_rand_val_run_x3_10_sva , psq_rand_val_run_x3_9_sva
      , psq_rand_val_run_x3_8_sva , psq_rand_val_run_x3_7_sva , psq_rand_val_run_x3_6_sva
      , psq_rand_val_run_x3_5_sva , psq_rand_val_run_x2_4_sva , psq_rand_val_run_x2_3_sva
      , psq_rand_val_run_x2_2_sva , psq_rand_val_run_x2_1_sva , psq_rand_val_run_x2_0_sva};
  assign psq_vecMul1_run_mul_cmp_3_b = {psq_run_py_not_2 , psq_rand_val2_run_x3_30_sva
      , psq_rand_val2_run_x3_29_sva , psq_rand_val2_run_x3_28_sva , psq_rand_val2_run_x3_27_sva
      , psq_rand_val2_run_x3_26_sva , psq_rand_val2_run_x3_25_sva , psq_rand_val2_run_x3_24_sva
      , psq_rand_val2_run_x3_23_sva , psq_rand_val2_run_x3_22_sva , psq_rand_val2_run_x3_21_sva
      , psq_rand_val2_run_x3_20_sva , psq_rand_val2_run_x3_19_sva , psq_rand_val2_run_x3_18_sva
      , psq_rand_val2_run_x3_17_sva , psq_rand_val2_run_x3_16_sva , psq_rand_val2_run_x3_15_sva
      , psq_rand_val2_run_x3_14_sva , psq_rand_val2_run_x3_13_sva , psq_rand_val2_run_x3_12_sva
      , psq_rand_val2_run_x3_11_sva , psq_rand_val2_run_x3_10_sva , psq_rand_val2_run_x3_9_sva
      , psq_rand_val2_run_x3_8_sva , psq_rand_val2_run_x3_7_sva , psq_rand_val2_run_x3_6_sva
      , psq_rand_val2_run_x3_5_sva , psq_rand_val2_run_x2_4_sva , psq_rand_val2_run_x2_3_sva
      , psq_rand_val2_run_x2_2_sva , psq_rand_val2_run_x2_1_sva , psq_rand_val2_run_x2_0_sva};
  assign psq_vecMul1_run_mul_cmp_2_b = {psq_run_px_not_3 , psq_rand_val_run_x3_30_sva
      , psq_rand_val_run_x3_29_sva , psq_rand_val_run_x3_28_sva , psq_rand_val_run_x3_27_sva
      , psq_rand_val_run_x3_26_sva , psq_rand_val_run_x3_25_sva , psq_rand_val_run_x3_24_sva
      , psq_rand_val_run_x3_23_sva , psq_rand_val_run_x3_22_sva , psq_rand_val_run_x3_21_sva
      , psq_rand_val_run_x3_20_sva , psq_rand_val_run_x3_19_sva , psq_rand_val_run_x3_18_sva
      , psq_rand_val_run_x3_17_sva , psq_rand_val_run_x3_16_sva , psq_rand_val_run_x3_15_sva
      , psq_rand_val_run_x3_14_sva , psq_rand_val_run_x3_13_sva , psq_rand_val_run_x3_12_sva
      , psq_rand_val_run_x3_11_sva , psq_rand_val_run_x3_10_sva , psq_rand_val_run_x3_9_sva
      , psq_rand_val_run_x3_8_sva , psq_rand_val_run_x3_7_sva , psq_rand_val_run_x3_6_sva
      , psq_rand_val_run_x3_5_sva , psq_rand_val_run_x2_4_sva , psq_rand_val_run_x2_3_sva
      , psq_rand_val_run_x2_2_sva , psq_rand_val_run_x2_1_sva , psq_rand_val_run_x2_0_sva};
  assign psq_vecMul1_run_mul_cmp_1_b = {psq_run_py_not_2 , psq_rand_val2_run_x3_30_sva
      , psq_rand_val2_run_x3_29_sva , psq_rand_val2_run_x3_28_sva , psq_rand_val2_run_x3_27_sva
      , psq_rand_val2_run_x3_26_sva , psq_rand_val2_run_x3_25_sva , psq_rand_val2_run_x3_24_sva
      , psq_rand_val2_run_x3_23_sva , psq_rand_val2_run_x3_22_sva , psq_rand_val2_run_x3_21_sva
      , psq_rand_val2_run_x3_20_sva , psq_rand_val2_run_x3_19_sva , psq_rand_val2_run_x3_18_sva
      , psq_rand_val2_run_x3_17_sva , psq_rand_val2_run_x3_16_sva , psq_rand_val2_run_x3_15_sva
      , psq_rand_val2_run_x3_14_sva , psq_rand_val2_run_x3_13_sva , psq_rand_val2_run_x3_12_sva
      , psq_rand_val2_run_x3_11_sva , psq_rand_val2_run_x3_10_sva , psq_rand_val2_run_x3_9_sva
      , psq_rand_val2_run_x3_8_sva , psq_rand_val2_run_x3_7_sva , psq_rand_val2_run_x3_6_sva
      , psq_rand_val2_run_x3_5_sva , psq_rand_val2_run_x2_4_sva , psq_rand_val2_run_x2_3_sva
      , psq_rand_val2_run_x2_2_sva , psq_rand_val2_run_x2_1_sva , psq_rand_val2_run_x2_0_sva};
  assign psq_vecMul1_run_mul_cmp_b = {psq_run_px_not_3 , psq_rand_val_run_x3_30_sva
      , psq_rand_val_run_x3_29_sva , psq_rand_val_run_x3_28_sva , psq_rand_val_run_x3_27_sva
      , psq_rand_val_run_x3_26_sva , psq_rand_val_run_x3_25_sva , psq_rand_val_run_x3_24_sva
      , psq_rand_val_run_x3_23_sva , psq_rand_val_run_x3_22_sva , psq_rand_val_run_x3_21_sva
      , psq_rand_val_run_x3_20_sva , psq_rand_val_run_x3_19_sva , psq_rand_val_run_x3_18_sva
      , psq_rand_val_run_x3_17_sva , psq_rand_val_run_x3_16_sva , psq_rand_val_run_x3_15_sva
      , psq_rand_val_run_x3_14_sva , psq_rand_val_run_x3_13_sva , psq_rand_val_run_x3_12_sva
      , psq_rand_val_run_x3_11_sva , psq_rand_val_run_x3_10_sva , psq_rand_val_run_x3_9_sva
      , psq_rand_val_run_x3_8_sva , psq_rand_val_run_x3_7_sva , psq_rand_val_run_x3_6_sva
      , psq_rand_val_run_x3_5_sva , psq_rand_val_run_x2_4_sva , psq_rand_val_run_x2_3_sva
      , psq_rand_val_run_x2_2_sva , psq_rand_val_run_x2_1_sva , psq_rand_val_run_x2_0_sva};
  assign rayOut_and_cse = run_wen & main_stage_0_4;
  assign and_itm = run_wen & main_stage_0_3;
  assign state2_and_cse = run_wen & (~ (fsm_output[0]));
  assign and_132_itm = run_wen & main_stage_0_2;
  assign nl_sampleAdd_run_acc_4_psp_sva_1 = deltAdd_run_acc_9_itm_2 + deltAdd_run_acc_8_itm_1;
  assign sampleAdd_run_acc_4_psp_sva_1 = nl_sampleAdd_run_acc_4_psp_sva_1[32:0];
  assign nl_sampleAdd_run_acc_3_psp_sva_1 = deltAdd_run_acc_7_itm_2 + deltAdd_run_acc_6_itm_1;
  assign sampleAdd_run_acc_3_psp_sva_1 = nl_sampleAdd_run_acc_3_psp_sva_1[32:0];
  assign nl_sampleAdd_run_acc_psp_sva_1 = deltAdd_run_acc_5_itm_2 + deltAdd_run_acc_itm_1;
  assign sampleAdd_run_acc_psp_sva_1 = nl_sampleAdd_run_acc_psp_sva_1[32:0];
  assign psq_rand_val2_run_x2_0_sva_4 = state2_0_sva ^ state2_17_sva ^ state2_4_sva;
  assign psq_rand_val2_run_x2_1_sva_4 = state2_1_sva ^ state2_18_sva ^ state2_5_sva;
  assign psq_rand_val2_run_x2_2_sva_4 = state2_2_sva ^ state2_19_sva ^ state2_6_sva;
  assign psq_rand_val2_run_x2_3_sva_4 = state2_3_sva ^ state2_20_sva ^ state2_7_sva;
  assign psq_rand_val2_run_x2_4_sva_4 = state2_4_sva ^ state2_21_sva ^ state2_8_sva;
  assign xor_cse = state2_5_sva ^ state2_22_sva ^ state2_9_sva;
  assign psq_rand_val2_run_x3_5_sva_4 = state2_0_sva ^ state2_17_sva ^ state2_4_sva
      ^ xor_cse;
  assign xor_cse_1 = state2_18_sva ^ state2_1_sva ^ state2_6_sva;
  assign psq_rand_val2_run_x3_6_sva_4 = state2_23_sva ^ state2_10_sva ^ state2_5_sva
      ^ xor_cse_1;
  assign xor_cse_2 = state2_11_sva ^ state2_24_sva ^ state2_7_sva;
  assign psq_rand_val2_run_x3_7_sva_4 = state2_2_sva ^ state2_19_sva ^ state2_6_sva
      ^ xor_cse_2;
  assign xor_cse_3 = state2_12_sva ^ state2_25_sva ^ state2_20_sva;
  assign psq_rand_val2_run_x3_8_sva_4 = state2_8_sva ^ state2_3_sva ^ state2_7_sva
      ^ xor_cse_3;
  assign xor_cse_4 = state2_13_sva ^ state2_26_sva ^ state2_9_sva;
  assign psq_rand_val2_run_x3_9_sva_4 = state2_4_sva ^ state2_21_sva ^ state2_8_sva
      ^ xor_cse_4;
  assign xor_cse_5 = state2_14_sva ^ state2_27_sva ^ state2_10_sva;
  assign psq_rand_val2_run_x3_10_sva_4 = xor_cse_5 ^ xor_cse;
  assign xor_cse_6 = state2_10_sva ^ state2_23_sva ^ state2_28_sva;
  assign psq_rand_val2_run_x3_11_sva_4 = state2_11_sva ^ state2_15_sva ^ state2_6_sva
      ^ xor_cse_6;
  assign xor_cse_7 = state2_16_sva ^ state2_29_sva ^ state2_12_sva;
  assign psq_rand_val2_run_x3_12_sva_4 = xor_cse_2 ^ xor_cse_7;
  assign xor_cse_8 = state2_17_sva ^ state2_0_sva ^ state2_13_sva ^ state2_30_sva;
  assign psq_rand_val2_run_x3_13_sva_4 = state2_8_sva ^ state2_25_sva ^ state2_12_sva
      ^ xor_cse_8;
  assign psq_rand_val2_run_x3_14_sva_4 = xor_cse_4 ^ state2_14_sva ^ state2_1_sva
      ^ state2_31_sva ^ state2_18_sva;
  assign psq_rand_val2_run_x3_15_sva_4 = state2_15_sva ^ state2_2_sva ^ xor_cse_5;
  assign psq_rand_val2_run_x3_16_sva_4 = state2_28_sva ^ state2_16_sva ^ state2_3_sva
      ^ state2_11_sva ^ state2_15_sva;
  assign psq_rand_val2_run_x3_17_sva_4 = state2_17_sva ^ state2_4_sva ^ xor_cse_7;
  assign psq_rand_val2_run_x3_18_sva_4 = state2_18_sva ^ state2_5_sva ^ xor_cse_8;
  assign psq_rand_val2_run_x3_19_sva_4 = state2_19_sva ^ state2_14_sva ^ state2_31_sva
      ^ xor_cse_1;
  assign psq_rand_val2_run_x3_20_sva_4 = state2_20_sva ^ state2_7_sva ^ state2_15_sva
      ^ state2_2_sva;
  assign psq_rand_val2_run_x3_21_sva_4 = state2_21_sva ^ state2_8_sva ^ state2_16_sva
      ^ state2_3_sva;
  assign psq_rand_val2_run_x3_22_sva_4 = state2_22_sva ^ state2_9_sva ^ state2_17_sva
      ^ state2_4_sva;
  assign psq_rand_val2_run_x3_23_sva_4 = state2_23_sva ^ state2_10_sva ^ state2_18_sva
      ^ state2_5_sva;
  assign psq_rand_val2_run_x3_24_sva_4 = state2_24_sva ^ state2_11_sva ^ state2_19_sva
      ^ state2_6_sva;
  assign psq_rand_val2_run_x3_25_sva_4 = state2_7_sva ^ xor_cse_3;
  assign psq_rand_val2_run_x3_26_sva_4 = state2_26_sva ^ state2_13_sva ^ state2_21_sva
      ^ state2_8_sva;
  assign psq_rand_val2_run_x3_27_sva_4 = state2_27_sva ^ state2_14_sva ^ state2_22_sva
      ^ state2_9_sva;
  assign psq_rand_val2_run_x3_28_sva_4 = state2_15_sva ^ xor_cse_6;
  assign psq_rand_val2_run_x3_29_sva_4 = state2_29_sva ^ state2_16_sva ^ state2_24_sva
      ^ state2_11_sva;
  assign psq_rand_val2_run_x3_30_sva_4 = state2_30_sva ^ state2_17_sva ^ state2_25_sva
      ^ state2_12_sva;
  assign psq_rand_val_run_x2_0_sva_4 = state1_0_sva ^ state1_17_sva ^ state1_4_sva;
  assign psq_rand_val_run_x2_1_sva_4 = state1_1_sva ^ state1_18_sva ^ state1_5_sva;
  assign psq_rand_val_run_x2_2_sva_4 = state1_2_sva ^ state1_19_sva ^ state1_6_sva;
  assign psq_rand_val_run_x2_3_sva_4 = state1_3_sva ^ state1_20_sva ^ state1_7_sva;
  assign psq_rand_val_run_x2_4_sva_4 = state1_4_sva ^ state1_21_sva ^ state1_8_sva;
  assign xor_cse_10 = state1_5_sva ^ state1_22_sva ^ state1_9_sva;
  assign psq_rand_val_run_x3_5_sva_4 = state1_0_sva ^ state1_17_sva ^ state1_4_sva
      ^ xor_cse_10;
  assign xor_cse_11 = state1_18_sva ^ state1_1_sva ^ state1_6_sva;
  assign psq_rand_val_run_x3_6_sva_4 = state1_23_sva ^ state1_10_sva ^ state1_5_sva
      ^ xor_cse_11;
  assign xor_cse_12 = state1_11_sva ^ state1_24_sva ^ state1_7_sva;
  assign psq_rand_val_run_x3_7_sva_4 = state1_2_sva ^ state1_19_sva ^ state1_6_sva
      ^ xor_cse_12;
  assign xor_cse_13 = state1_12_sva ^ state1_25_sva ^ state1_20_sva;
  assign psq_rand_val_run_x3_8_sva_4 = state1_8_sva ^ state1_3_sva ^ state1_7_sva
      ^ xor_cse_13;
  assign xor_cse_14 = state1_13_sva ^ state1_26_sva ^ state1_9_sva;
  assign psq_rand_val_run_x3_9_sva_4 = state1_4_sva ^ state1_21_sva ^ state1_8_sva
      ^ xor_cse_14;
  assign xor_cse_15 = state1_14_sva ^ state1_27_sva ^ state1_10_sva;
  assign psq_rand_val_run_x3_10_sva_4 = xor_cse_15 ^ xor_cse_10;
  assign xor_cse_16 = state1_10_sva ^ state1_23_sva ^ state1_28_sva;
  assign psq_rand_val_run_x3_11_sva_4 = state1_11_sva ^ state1_15_sva ^ state1_6_sva
      ^ xor_cse_16;
  assign xor_cse_17 = state1_16_sva ^ state1_29_sva ^ state1_12_sva;
  assign psq_rand_val_run_x3_12_sva_4 = xor_cse_12 ^ xor_cse_17;
  assign xor_cse_18 = state1_17_sva ^ state1_0_sva ^ state1_13_sva ^ state1_30_sva;
  assign psq_rand_val_run_x3_13_sva_4 = state1_8_sva ^ state1_25_sva ^ state1_12_sva
      ^ xor_cse_18;
  assign psq_rand_val_run_x3_14_sva_4 = xor_cse_14 ^ state1_14_sva ^ state1_1_sva
      ^ state1_31_sva ^ state1_18_sva;
  assign psq_rand_val_run_x3_15_sva_4 = state1_15_sva ^ state1_2_sva ^ xor_cse_15;
  assign psq_rand_val_run_x3_16_sva_4 = state1_28_sva ^ state1_16_sva ^ state1_3_sva
      ^ state1_11_sva ^ state1_15_sva;
  assign psq_rand_val_run_x3_17_sva_4 = state1_17_sva ^ state1_4_sva ^ xor_cse_17;
  assign psq_rand_val_run_x3_18_sva_4 = state1_18_sva ^ state1_5_sva ^ xor_cse_18;
  assign psq_rand_val_run_x3_19_sva_4 = state1_19_sva ^ state1_14_sva ^ state1_31_sva
      ^ xor_cse_11;
  assign psq_rand_val_run_x3_20_sva_4 = state1_20_sva ^ state1_7_sva ^ state1_15_sva
      ^ state1_2_sva;
  assign psq_rand_val_run_x3_21_sva_4 = state1_21_sva ^ state1_8_sva ^ state1_16_sva
      ^ state1_3_sva;
  assign psq_rand_val_run_x3_22_sva_4 = state1_22_sva ^ state1_9_sva ^ state1_17_sva
      ^ state1_4_sva;
  assign psq_rand_val_run_x3_23_sva_4 = state1_23_sva ^ state1_10_sva ^ state1_18_sva
      ^ state1_5_sva;
  assign psq_rand_val_run_x3_24_sva_4 = state1_24_sva ^ state1_11_sva ^ state1_19_sva
      ^ state1_6_sva;
  assign psq_rand_val_run_x3_25_sva_4 = state1_7_sva ^ xor_cse_13;
  assign psq_rand_val_run_x3_26_sva_4 = state1_26_sva ^ state1_13_sva ^ state1_21_sva
      ^ state1_8_sva;
  assign psq_rand_val_run_x3_27_sva_4 = state1_27_sva ^ state1_14_sva ^ state1_22_sva
      ^ state1_9_sva;
  assign psq_rand_val_run_x3_28_sva_4 = state1_15_sva ^ xor_cse_16;
  assign psq_rand_val_run_x3_29_sva_4 = state1_29_sva ^ state1_16_sva ^ state1_24_sva
      ^ state1_11_sva;
  assign psq_rand_val_run_x3_30_sva_4 = state1_30_sva ^ state1_17_sva ^ state1_25_sva
      ^ state1_12_sva;
  assign xor_cse_20 = state2_18_sva ^ state2_31_sva ^ state2_26_sva;
  assign xor_cse_21 = state1_18_sva ^ state1_31_sva ^ state1_26_sva;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayOut_rsci_idat_20_10 <= 11'b00000000000;
      rayOut_rsci_idat_41_31 <= 11'b00000000000;
      rayOut_rsci_idat_62_52 <= 11'b00000000000;
      rayOut_rsci_idat_85_64 <= 22'b0000000000000000000000;
      rayOut_rsci_idat_96_86 <= 11'b00000000000;
      rayOut_rsci_idat_119_98 <= 22'b0000000000000000000000;
      rayOut_rsci_idat_130_120 <= 11'b00000000000;
      rayOut_rsci_idat_153_132 <= 22'b0000000000000000000000;
      rayOut_rsci_idat_164_154 <= 11'b00000000000;
      paramsOut_rsci_idat_10_0 <= 11'b00000000000;
      paramsOut_rsci_idat_91_11 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      paramsOut_rsci_idat_92 <= 1'b0;
    end
    else if ( rayOut_and_cse ) begin
      rayOut_rsci_idat_20_10 <= paramsIn_crt_sva_3_170_138[10:0];
      rayOut_rsci_idat_41_31 <= paramsIn_crt_sva_3_170_138[21:11];
      rayOut_rsci_idat_62_52 <= paramsIn_crt_sva_3_170_138[32:22];
      rayOut_rsci_idat_85_64 <= sampleAdd_run_acc_psp_sva_1[21:0];
      rayOut_rsci_idat_96_86 <= nl_rayOut_rsci_idat_96_86[10:0];
      rayOut_rsci_idat_119_98 <= sampleAdd_run_acc_3_psp_sva_1[21:0];
      rayOut_rsci_idat_130_120 <= nl_rayOut_rsci_idat_130_120[10:0];
      rayOut_rsci_idat_153_132 <= sampleAdd_run_acc_4_psp_sva_1[21:0];
      rayOut_rsci_idat_164_154 <= nl_rayOut_rsci_idat_164_154[10:0];
      paramsOut_rsci_idat_10_0 <= paramsIn_crt_sva_3_10_0;
      paramsOut_rsci_idat_91_11 <= paramsIn_crt_sva_3_93_13;
      paramsOut_rsci_idat_92 <= loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_rayOut_rsci_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      psq_rand_val2_run_x2_0_sva <= 1'b0;
      psq_rand_val2_run_x2_1_sva <= 1'b0;
      psq_rand_val2_run_x2_2_sva <= 1'b0;
      psq_rand_val2_run_x2_3_sva <= 1'b0;
      psq_rand_val2_run_x2_4_sva <= 1'b0;
      psq_rand_val2_run_x3_5_sva <= 1'b0;
      psq_rand_val2_run_x3_6_sva <= 1'b0;
      psq_rand_val2_run_x3_7_sva <= 1'b0;
      psq_rand_val2_run_x3_8_sva <= 1'b0;
      psq_rand_val2_run_x3_9_sva <= 1'b0;
      psq_rand_val2_run_x3_10_sva <= 1'b0;
      psq_rand_val2_run_x3_11_sva <= 1'b0;
      psq_rand_val2_run_x3_12_sva <= 1'b0;
      psq_rand_val2_run_x3_13_sva <= 1'b0;
      psq_rand_val2_run_x3_14_sva <= 1'b0;
      psq_rand_val2_run_x3_15_sva <= 1'b0;
      psq_rand_val2_run_x3_16_sva <= 1'b0;
      psq_rand_val2_run_x3_17_sva <= 1'b0;
      psq_rand_val2_run_x3_18_sva <= 1'b0;
      psq_rand_val2_run_x3_19_sva <= 1'b0;
      psq_rand_val2_run_x3_20_sva <= 1'b0;
      psq_rand_val2_run_x3_21_sva <= 1'b0;
      psq_rand_val2_run_x3_22_sva <= 1'b0;
      psq_rand_val2_run_x3_23_sva <= 1'b0;
      psq_rand_val2_run_x3_24_sva <= 1'b0;
      psq_rand_val2_run_x3_25_sva <= 1'b0;
      psq_rand_val2_run_x3_26_sva <= 1'b0;
      psq_rand_val2_run_x3_27_sva <= 1'b0;
      psq_rand_val2_run_x3_28_sva <= 1'b0;
      psq_rand_val2_run_x3_29_sva <= 1'b0;
      psq_rand_val2_run_x3_30_sva <= 1'b0;
      psq_run_py_not_2 <= 1'b0;
      psq_vecMul1_run_mul_cmp_5_a <= 25'b0000000000000000000000000;
      psq_rand_val_run_x2_0_sva <= 1'b0;
      psq_rand_val_run_x2_1_sva <= 1'b0;
      psq_rand_val_run_x2_2_sva <= 1'b0;
      psq_rand_val_run_x2_3_sva <= 1'b0;
      psq_rand_val_run_x2_4_sva <= 1'b0;
      psq_rand_val_run_x3_5_sva <= 1'b0;
      psq_rand_val_run_x3_6_sva <= 1'b0;
      psq_rand_val_run_x3_7_sva <= 1'b0;
      psq_rand_val_run_x3_8_sva <= 1'b0;
      psq_rand_val_run_x3_9_sva <= 1'b0;
      psq_rand_val_run_x3_10_sva <= 1'b0;
      psq_rand_val_run_x3_11_sva <= 1'b0;
      psq_rand_val_run_x3_12_sva <= 1'b0;
      psq_rand_val_run_x3_13_sva <= 1'b0;
      psq_rand_val_run_x3_14_sva <= 1'b0;
      psq_rand_val_run_x3_15_sva <= 1'b0;
      psq_rand_val_run_x3_16_sva <= 1'b0;
      psq_rand_val_run_x3_17_sva <= 1'b0;
      psq_rand_val_run_x3_18_sva <= 1'b0;
      psq_rand_val_run_x3_19_sva <= 1'b0;
      psq_rand_val_run_x3_20_sva <= 1'b0;
      psq_rand_val_run_x3_21_sva <= 1'b0;
      psq_rand_val_run_x3_22_sva <= 1'b0;
      psq_rand_val_run_x3_23_sva <= 1'b0;
      psq_rand_val_run_x3_24_sva <= 1'b0;
      psq_rand_val_run_x3_25_sva <= 1'b0;
      psq_rand_val_run_x3_26_sva <= 1'b0;
      psq_rand_val_run_x3_27_sva <= 1'b0;
      psq_rand_val_run_x3_28_sva <= 1'b0;
      psq_rand_val_run_x3_29_sva <= 1'b0;
      psq_rand_val_run_x3_30_sva <= 1'b0;
      psq_run_px_not_3 <= 1'b0;
      psq_vecMul1_run_mul_cmp_4_a <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_3_a <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_2_a <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_1_a <= 25'b0000000000000000000000000;
      psq_vecMul1_run_mul_cmp_a <= 25'b0000000000000000000000000;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      deltUMul_run_mul_2_itm_1 <= 33'b000000000000000000000000000000000;
      deltVMul_run_mul_2_itm_1 <= 33'b000000000000000000000000000000000;
      deltUMul_run_mul_1_itm_1 <= 33'b000000000000000000000000000000000;
      deltVMul_run_mul_1_itm_1 <= 33'b000000000000000000000000000000000;
      deltUMul_run_mul_itm_1 <= 33'b000000000000000000000000000000000;
      deltVMul_run_mul_itm_1 <= 33'b000000000000000000000000000000000;
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_1 <= 1'b0;
      paramsIn_crt_sva_1_269_138 <= 132'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      paramsIn_crt_sva_1_10_0 <= 11'b00000000000;
      paramsIn_crt_sva_1_93_13 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_rayOut_rsci_ivld_run_psct_cse <= main_stage_0_4;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b1;
      psq_rand_val2_run_x2_0_sva <= psq_rand_val2_run_x2_0_sva_4;
      psq_rand_val2_run_x2_1_sva <= psq_rand_val2_run_x2_1_sva_4;
      psq_rand_val2_run_x2_2_sva <= psq_rand_val2_run_x2_2_sva_4;
      psq_rand_val2_run_x2_3_sva <= psq_rand_val2_run_x2_3_sva_4;
      psq_rand_val2_run_x2_4_sva <= psq_rand_val2_run_x2_4_sva_4;
      psq_rand_val2_run_x3_5_sva <= psq_rand_val2_run_x3_5_sva_4;
      psq_rand_val2_run_x3_6_sva <= psq_rand_val2_run_x3_6_sva_4;
      psq_rand_val2_run_x3_7_sva <= psq_rand_val2_run_x3_7_sva_4;
      psq_rand_val2_run_x3_8_sva <= psq_rand_val2_run_x3_8_sva_4;
      psq_rand_val2_run_x3_9_sva <= psq_rand_val2_run_x3_9_sva_4;
      psq_rand_val2_run_x3_10_sva <= psq_rand_val2_run_x3_10_sva_4;
      psq_rand_val2_run_x3_11_sva <= psq_rand_val2_run_x3_11_sva_4;
      psq_rand_val2_run_x3_12_sva <= psq_rand_val2_run_x3_12_sva_4;
      psq_rand_val2_run_x3_13_sva <= psq_rand_val2_run_x3_13_sva_4;
      psq_rand_val2_run_x3_14_sva <= psq_rand_val2_run_x3_14_sva_4;
      psq_rand_val2_run_x3_15_sva <= psq_rand_val2_run_x3_15_sva_4;
      psq_rand_val2_run_x3_16_sva <= psq_rand_val2_run_x3_16_sva_4;
      psq_rand_val2_run_x3_17_sva <= psq_rand_val2_run_x3_17_sva_4;
      psq_rand_val2_run_x3_18_sva <= psq_rand_val2_run_x3_18_sva_4;
      psq_rand_val2_run_x3_19_sva <= psq_rand_val2_run_x3_19_sva_4;
      psq_rand_val2_run_x3_20_sva <= psq_rand_val2_run_x3_20_sva_4;
      psq_rand_val2_run_x3_21_sva <= psq_rand_val2_run_x3_21_sva_4;
      psq_rand_val2_run_x3_22_sva <= psq_rand_val2_run_x3_22_sva_4;
      psq_rand_val2_run_x3_23_sva <= psq_rand_val2_run_x3_23_sva_4;
      psq_rand_val2_run_x3_24_sva <= psq_rand_val2_run_x3_24_sva_4;
      psq_rand_val2_run_x3_25_sva <= psq_rand_val2_run_x3_25_sva_4;
      psq_rand_val2_run_x3_26_sva <= psq_rand_val2_run_x3_26_sva_4;
      psq_rand_val2_run_x3_27_sva <= psq_rand_val2_run_x3_27_sva_4;
      psq_rand_val2_run_x3_28_sva <= psq_rand_val2_run_x3_28_sva_4;
      psq_rand_val2_run_x3_29_sva <= psq_rand_val2_run_x3_29_sva_4;
      psq_rand_val2_run_x3_30_sva <= psq_rand_val2_run_x3_30_sva_4;
      psq_run_py_not_2 <= ~(state2_13_sva ^ xor_cse_20);
      psq_vecMul1_run_mul_cmp_5_a <= paramsIn_rsci_idat_mxwt[323:299];
      psq_rand_val_run_x2_0_sva <= psq_rand_val_run_x2_0_sva_4;
      psq_rand_val_run_x2_1_sva <= psq_rand_val_run_x2_1_sva_4;
      psq_rand_val_run_x2_2_sva <= psq_rand_val_run_x2_2_sva_4;
      psq_rand_val_run_x2_3_sva <= psq_rand_val_run_x2_3_sva_4;
      psq_rand_val_run_x2_4_sva <= psq_rand_val_run_x2_4_sva_4;
      psq_rand_val_run_x3_5_sva <= psq_rand_val_run_x3_5_sva_4;
      psq_rand_val_run_x3_6_sva <= psq_rand_val_run_x3_6_sva_4;
      psq_rand_val_run_x3_7_sva <= psq_rand_val_run_x3_7_sva_4;
      psq_rand_val_run_x3_8_sva <= psq_rand_val_run_x3_8_sva_4;
      psq_rand_val_run_x3_9_sva <= psq_rand_val_run_x3_9_sva_4;
      psq_rand_val_run_x3_10_sva <= psq_rand_val_run_x3_10_sva_4;
      psq_rand_val_run_x3_11_sva <= psq_rand_val_run_x3_11_sva_4;
      psq_rand_val_run_x3_12_sva <= psq_rand_val_run_x3_12_sva_4;
      psq_rand_val_run_x3_13_sva <= psq_rand_val_run_x3_13_sva_4;
      psq_rand_val_run_x3_14_sva <= psq_rand_val_run_x3_14_sva_4;
      psq_rand_val_run_x3_15_sva <= psq_rand_val_run_x3_15_sva_4;
      psq_rand_val_run_x3_16_sva <= psq_rand_val_run_x3_16_sva_4;
      psq_rand_val_run_x3_17_sva <= psq_rand_val_run_x3_17_sva_4;
      psq_rand_val_run_x3_18_sva <= psq_rand_val_run_x3_18_sva_4;
      psq_rand_val_run_x3_19_sva <= psq_rand_val_run_x3_19_sva_4;
      psq_rand_val_run_x3_20_sva <= psq_rand_val_run_x3_20_sva_4;
      psq_rand_val_run_x3_21_sva <= psq_rand_val_run_x3_21_sva_4;
      psq_rand_val_run_x3_22_sva <= psq_rand_val_run_x3_22_sva_4;
      psq_rand_val_run_x3_23_sva <= psq_rand_val_run_x3_23_sva_4;
      psq_rand_val_run_x3_24_sva <= psq_rand_val_run_x3_24_sva_4;
      psq_rand_val_run_x3_25_sva <= psq_rand_val_run_x3_25_sva_4;
      psq_rand_val_run_x3_26_sva <= psq_rand_val_run_x3_26_sva_4;
      psq_rand_val_run_x3_27_sva <= psq_rand_val_run_x3_27_sva_4;
      psq_rand_val_run_x3_28_sva <= psq_rand_val_run_x3_28_sva_4;
      psq_rand_val_run_x3_29_sva <= psq_rand_val_run_x3_29_sva_4;
      psq_rand_val_run_x3_30_sva <= psq_rand_val_run_x3_30_sva_4;
      psq_run_px_not_3 <= ~(state1_13_sva ^ xor_cse_21);
      psq_vecMul1_run_mul_cmp_4_a <= paramsIn_rsci_idat_mxwt[273:249];
      psq_vecMul1_run_mul_cmp_3_a <= paramsIn_rsci_idat_mxwt[348:324];
      psq_vecMul1_run_mul_cmp_2_a <= paramsIn_rsci_idat_mxwt[298:274];
      psq_vecMul1_run_mul_cmp_1_a <= paramsIn_rsci_idat_mxwt[373:349];
      psq_vecMul1_run_mul_cmp_a <= paramsIn_rsci_idat_mxwt[248:224];
      main_stage_0_2 <= fsm_output[1];
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      deltUMul_run_mul_2_itm_1 <= nl_deltUMul_run_mul_2_itm_1[32:0];
      deltVMul_run_mul_2_itm_1 <= nl_deltVMul_run_mul_2_itm_1[32:0];
      deltUMul_run_mul_1_itm_1 <= nl_deltUMul_run_mul_1_itm_1[32:0];
      deltVMul_run_mul_1_itm_1 <= nl_deltVMul_run_mul_1_itm_1[32:0];
      deltUMul_run_mul_itm_1 <= nl_deltUMul_run_mul_itm_1[32:0];
      deltVMul_run_mul_itm_1 <= nl_deltVMul_run_mul_itm_1[32:0];
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_1 <= loopIndicesIn_rsci_idat_mxwt[22];
      paramsIn_crt_sva_1_269_138 <= paramsIn_rsci_idat_mxwt[223:92];
      paramsIn_crt_sva_1_10_0 <= paramsIn_rsci_idat_mxwt[10:0];
      paramsIn_crt_sva_1_93_13 <= paramsIn_rsci_idat_mxwt[91:11];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_sva_3_170_138 <= 33'b000000000000000000000000000000000;
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_3 <= 1'b0;
      paramsIn_crt_sva_3_10_0 <= 11'b00000000000;
      paramsIn_crt_sva_3_93_13 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      deltAdd_run_acc_9_itm_2 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_8_itm_1 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_7_itm_2 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_6_itm_1 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_5_itm_2 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_itm_1 <= 33'b000000000000000000000000000000000;
    end
    else if ( and_itm ) begin
      paramsIn_crt_sva_3_170_138 <= paramsIn_crt_sva_2_269_138[32:0];
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_3 <= loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_2;
      paramsIn_crt_sva_3_10_0 <= paramsIn_crt_sva_2_10_0;
      paramsIn_crt_sva_3_93_13 <= paramsIn_crt_sva_2_93_13;
      deltAdd_run_acc_9_itm_2 <= deltAdd_run_acc_9_itm_1;
      deltAdd_run_acc_8_itm_1 <= nl_deltAdd_run_acc_8_itm_1[32:0];
      deltAdd_run_acc_7_itm_2 <= deltAdd_run_acc_7_itm_1;
      deltAdd_run_acc_6_itm_1 <= nl_deltAdd_run_acc_6_itm_1[32:0];
      deltAdd_run_acc_5_itm_2 <= deltAdd_run_acc_5_itm_1;
      deltAdd_run_acc_itm_1 <= nl_deltAdd_run_acc_itm_1[32:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state2_0_sva <= 1'b0;
      state2_1_sva <= 1'b0;
      state2_2_sva <= 1'b0;
      state2_3_sva <= 1'b0;
      state2_4_sva <= 1'b1;
      state2_5_sva <= 1'b0;
      state2_6_sva <= 1'b0;
      state2_7_sva <= 1'b1;
      state2_8_sva <= 1'b0;
      state2_9_sva <= 1'b0;
      state2_10_sva <= 1'b1;
      state2_11_sva <= 1'b1;
      state2_12_sva <= 1'b0;
      state2_13_sva <= 1'b1;
      state2_14_sva <= 1'b1;
      state2_16_sva <= 1'b0;
      state2_15_sva <= 1'b1;
      state2_31_sva <= 1'b0;
      state2_18_sva <= 1'b1;
      state2_30_sva <= 1'b0;
      state2_17_sva <= 1'b1;
      state2_29_sva <= 1'b0;
      state2_28_sva <= 1'b0;
      state2_27_sva <= 1'b0;
      state2_26_sva <= 1'b0;
      state2_25_sva <= 1'b1;
      state2_24_sva <= 1'b0;
      state2_23_sva <= 1'b0;
      state2_22_sva <= 1'b1;
      state2_21_sva <= 1'b0;
      state2_20_sva <= 1'b1;
      state2_19_sva <= 1'b0;
      state1_0_sva <= 1'b1;
      state1_1_sva <= 1'b0;
      state1_2_sva <= 1'b1;
      state1_3_sva <= 1'b1;
      state1_4_sva <= 1'b0;
      state1_5_sva <= 1'b0;
      state1_6_sva <= 1'b0;
      state1_7_sva <= 1'b0;
      state1_8_sva <= 1'b0;
      state1_9_sva <= 1'b0;
      state1_10_sva <= 1'b1;
      state1_11_sva <= 1'b1;
      state1_12_sva <= 1'b1;
      state1_13_sva <= 1'b1;
      state1_14_sva <= 1'b0;
      state1_16_sva <= 1'b1;
      state1_15_sva <= 1'b1;
      state1_31_sva <= 1'b0;
      state1_18_sva <= 1'b1;
      state1_30_sva <= 1'b0;
      state1_17_sva <= 1'b0;
      state1_29_sva <= 1'b0;
      state1_28_sva <= 1'b0;
      state1_27_sva <= 1'b0;
      state1_26_sva <= 1'b0;
      state1_25_sva <= 1'b0;
      state1_24_sva <= 1'b0;
      state1_23_sva <= 1'b0;
      state1_22_sva <= 1'b0;
      state1_21_sva <= 1'b0;
      state1_20_sva <= 1'b0;
      state1_19_sva <= 1'b0;
    end
    else if ( state2_and_cse ) begin
      state2_0_sva <= psq_rand_val2_run_x2_0_sva_4;
      state2_1_sva <= psq_rand_val2_run_x2_1_sva_4;
      state2_2_sva <= psq_rand_val2_run_x2_2_sva_4;
      state2_3_sva <= psq_rand_val2_run_x2_3_sva_4;
      state2_4_sva <= psq_rand_val2_run_x2_4_sva_4;
      state2_5_sva <= psq_rand_val2_run_x3_5_sva_4;
      state2_6_sva <= psq_rand_val2_run_x3_6_sva_4;
      state2_7_sva <= psq_rand_val2_run_x3_7_sva_4;
      state2_8_sva <= psq_rand_val2_run_x3_8_sva_4;
      state2_9_sva <= psq_rand_val2_run_x3_9_sva_4;
      state2_10_sva <= psq_rand_val2_run_x3_10_sva_4;
      state2_11_sva <= psq_rand_val2_run_x3_11_sva_4;
      state2_12_sva <= psq_rand_val2_run_x3_12_sva_4;
      state2_13_sva <= psq_rand_val2_run_x3_13_sva_4;
      state2_14_sva <= psq_rand_val2_run_x3_14_sva_4;
      state2_16_sva <= psq_rand_val2_run_x3_16_sva_4;
      state2_15_sva <= psq_rand_val2_run_x3_15_sva_4;
      state2_31_sva <= state2_13_sva ^ xor_cse_20;
      state2_18_sva <= psq_rand_val2_run_x3_18_sva_4;
      state2_30_sva <= psq_rand_val2_run_x3_30_sva_4;
      state2_17_sva <= psq_rand_val2_run_x3_17_sva_4;
      state2_29_sva <= psq_rand_val2_run_x3_29_sva_4;
      state2_28_sva <= psq_rand_val2_run_x3_28_sva_4;
      state2_27_sva <= psq_rand_val2_run_x3_27_sva_4;
      state2_26_sva <= psq_rand_val2_run_x3_26_sva_4;
      state2_25_sva <= psq_rand_val2_run_x3_25_sva_4;
      state2_24_sva <= psq_rand_val2_run_x3_24_sva_4;
      state2_23_sva <= psq_rand_val2_run_x3_23_sva_4;
      state2_22_sva <= psq_rand_val2_run_x3_22_sva_4;
      state2_21_sva <= psq_rand_val2_run_x3_21_sva_4;
      state2_20_sva <= psq_rand_val2_run_x3_20_sva_4;
      state2_19_sva <= psq_rand_val2_run_x3_19_sva_4;
      state1_0_sva <= psq_rand_val_run_x2_0_sva_4;
      state1_1_sva <= psq_rand_val_run_x2_1_sva_4;
      state1_2_sva <= psq_rand_val_run_x2_2_sva_4;
      state1_3_sva <= psq_rand_val_run_x2_3_sva_4;
      state1_4_sva <= psq_rand_val_run_x2_4_sva_4;
      state1_5_sva <= psq_rand_val_run_x3_5_sva_4;
      state1_6_sva <= psq_rand_val_run_x3_6_sva_4;
      state1_7_sva <= psq_rand_val_run_x3_7_sva_4;
      state1_8_sva <= psq_rand_val_run_x3_8_sva_4;
      state1_9_sva <= psq_rand_val_run_x3_9_sva_4;
      state1_10_sva <= psq_rand_val_run_x3_10_sva_4;
      state1_11_sva <= psq_rand_val_run_x3_11_sva_4;
      state1_12_sva <= psq_rand_val_run_x3_12_sva_4;
      state1_13_sva <= psq_rand_val_run_x3_13_sva_4;
      state1_14_sva <= psq_rand_val_run_x3_14_sva_4;
      state1_16_sva <= psq_rand_val_run_x3_16_sva_4;
      state1_15_sva <= psq_rand_val_run_x3_15_sva_4;
      state1_31_sva <= state1_13_sva ^ xor_cse_21;
      state1_18_sva <= psq_rand_val_run_x3_18_sva_4;
      state1_30_sva <= psq_rand_val_run_x3_30_sva_4;
      state1_17_sva <= psq_rand_val_run_x3_17_sva_4;
      state1_29_sva <= psq_rand_val_run_x3_29_sva_4;
      state1_28_sva <= psq_rand_val_run_x3_28_sva_4;
      state1_27_sva <= psq_rand_val_run_x3_27_sva_4;
      state1_26_sva <= psq_rand_val_run_x3_26_sva_4;
      state1_25_sva <= psq_rand_val_run_x3_25_sva_4;
      state1_24_sva <= psq_rand_val_run_x3_24_sva_4;
      state1_23_sva <= psq_rand_val_run_x3_23_sva_4;
      state1_22_sva <= psq_rand_val_run_x3_22_sva_4;
      state1_21_sva <= psq_rand_val_run_x3_21_sva_4;
      state1_20_sva <= psq_rand_val_run_x3_20_sva_4;
      state1_19_sva <= psq_rand_val_run_x3_19_sva_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      paramsIn_crt_sva_2_269_138 <= 132'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_2 <= 1'b0;
      deltAdd_run_acc_9_itm_1 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_7_itm_1 <= 33'b000000000000000000000000000000000;
      deltAdd_run_acc_5_itm_1 <= 33'b000000000000000000000000000000000;
      paramsIn_crt_sva_2_10_0 <= 11'b00000000000;
      paramsIn_crt_sva_2_93_13 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_132_itm ) begin
      paramsIn_crt_sva_2_269_138 <= paramsIn_crt_sva_1_269_138;
      loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_2 <= loopIndicesIn_lastsamp_slc_loopIndicesIn_crt_22_itm_1;
      deltAdd_run_acc_9_itm_1 <= nl_deltAdd_run_acc_9_itm_1[32:0];
      deltAdd_run_acc_7_itm_1 <= nl_deltAdd_run_acc_7_itm_1[32:0];
      deltAdd_run_acc_5_itm_1 <= nl_deltAdd_run_acc_5_itm_1[32:0];
      paramsIn_crt_sva_2_10_0 <= paramsIn_crt_sva_1_10_0;
      paramsIn_crt_sva_2_93_13 <= paramsIn_crt_sva_1_93_13;
    end
  end
  assign nl_rayOut_rsci_idat_96_86  = (sampleAdd_run_acc_psp_sva_1[32:22]) - (paramsIn_crt_sva_3_170_138[10:0]);
  assign nl_rayOut_rsci_idat_130_120  = (sampleAdd_run_acc_3_psp_sva_1[32:22]) -
      (paramsIn_crt_sva_3_170_138[21:11]);
  assign nl_rayOut_rsci_idat_164_154  = (sampleAdd_run_acc_4_psp_sva_1[32:22]) -
      (paramsIn_crt_sva_3_170_138[32:22]);
  assign nl_deltUMul_run_mul_2_itm_1  = $signed((paramsIn_rsci_idat_mxwt[298:274]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[10:0]));
  assign nl_deltVMul_run_mul_2_itm_1  = $signed((paramsIn_rsci_idat_mxwt[373:349]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[21:11]));
  assign nl_deltUMul_run_mul_1_itm_1  = $signed((paramsIn_rsci_idat_mxwt[273:249]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[10:0]));
  assign nl_deltVMul_run_mul_1_itm_1  = $signed((paramsIn_rsci_idat_mxwt[348:324]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[21:11]));
  assign nl_deltUMul_run_mul_itm_1  = $signed((paramsIn_rsci_idat_mxwt[248:224]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[10:0]));
  assign nl_deltVMul_run_mul_itm_1  = $signed((paramsIn_rsci_idat_mxwt[323:299]))
      * $signed(conv_u2s_11_12(loopIndicesIn_rsci_idat_mxwt[21:11]));
  assign nl_psq_run_acc_2_nl = psq_vecMul1_run_mul_cmp_2_z_oreg + psq_vecMul1_run_mul_cmp_1_z_oreg;
  assign psq_run_acc_2_nl = nl_psq_run_acc_2_nl[24:0];
  assign nl_deltAdd_run_acc_8_itm_1  = (paramsIn_crt_sva_2_269_138[131:99]) + conv_s2s_25_33(psq_run_acc_2_nl);
  assign nl_psq_run_acc_1_nl = psq_vecMul1_run_mul_cmp_4_z_oreg + psq_vecMul1_run_mul_cmp_3_z_oreg;
  assign psq_run_acc_1_nl = nl_psq_run_acc_1_nl[24:0];
  assign nl_deltAdd_run_acc_6_itm_1  = (paramsIn_crt_sva_2_269_138[98:66]) + conv_s2s_25_33(psq_run_acc_1_nl);
  assign nl_psq_run_acc_nl = psq_vecMul1_run_mul_cmp_z_oreg + psq_vecMul1_run_mul_cmp_5_z_oreg;
  assign psq_run_acc_nl = nl_psq_run_acc_nl[24:0];
  assign nl_deltAdd_run_acc_itm_1  = (paramsIn_crt_sva_2_269_138[65:33]) + conv_s2s_25_33(psq_run_acc_nl);
  assign nl_deltAdd_run_acc_9_itm_1  = deltUMul_run_mul_2_itm_1 + deltVMul_run_mul_2_itm_1;
  assign nl_deltAdd_run_acc_7_itm_1  = deltUMul_run_mul_1_itm_1 + deltVMul_run_mul_1_itm_1;
  assign nl_deltAdd_run_acc_5_itm_1  = deltUMul_run_mul_itm_1 + deltVMul_run_mul_itm_1;

  function automatic [32:0] conv_s2s_25_33 ;
    input [24:0]  vector ;
  begin
    conv_s2s_25_33 = {{8{vector[24]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib_run
// ------------------------------------------------------------------


module LoopDistrib_run (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy,
      attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld, accumalated_color_chan_in_rsc_rdy,
      attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      ray_out_loopone_rsc_dat, ray_out_loopone_rsc_vld, ray_out_loopone_rsc_rdy,
      ray_out_looptwo_rsc_dat, ray_out_looptwo_rsc_vld, ray_out_looptwo_rsc_rdy,
      ray_out_worldhit_rsc_dat, ray_out_worldhit_rsc_vld, ray_out_worldhit_rsc_rdy,
      quad_out_loopone_rsc_dat, quad_out_loopone_rsc_vld, quad_out_loopone_rsc_rdy,
      quad_out_looptwo_rsc_dat, quad_out_looptwo_rsc_vld, quad_out_looptwo_rsc_rdy,
      quad_max_outone_rsc_dat, quad_max_outone_rsc_vld, quad_max_outone_rsc_rdy,
      quad_max_outtwo_rsc_dat, quad_max_outtwo_rsc_vld, quad_max_outtwo_rsc_rdy,
      params_out_rsc_dat, params_out_rsc_vld, params_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [165:0] ray_out_loopone_rsc_dat;
  output ray_out_loopone_rsc_vld;
  input ray_out_loopone_rsc_rdy;
  output [165:0] ray_out_looptwo_rsc_dat;
  output ray_out_looptwo_rsc_vld;
  input ray_out_looptwo_rsc_rdy;
  output [165:0] ray_out_worldhit_rsc_dat;
  output ray_out_worldhit_rsc_vld;
  input ray_out_worldhit_rsc_rdy;
  output [376:0] quad_out_loopone_rsc_dat;
  output quad_out_loopone_rsc_vld;
  input quad_out_loopone_rsc_rdy;
  output [376:0] quad_out_looptwo_rsc_dat;
  output quad_out_looptwo_rsc_vld;
  input quad_out_looptwo_rsc_rdy;
  output [10:0] quad_max_outone_rsc_dat;
  output quad_max_outone_rsc_vld;
  input quad_max_outone_rsc_rdy;
  output [10:0] quad_max_outtwo_rsc_dat;
  output quad_max_outtwo_rsc_vld;
  input quad_max_outtwo_rsc_rdy;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire ray_in_rsci_wen_comp;
  wire [165:0] ray_in_rsci_idat_mxwt;
  wire params_in_rsci_wen_comp;
  wire [92:0] params_in_rsci_idat_mxwt;
  wire quads_rsci_wen_comp;
  wire [376:0] quads_rsci_idat_mxwt;
  wire attenuation_chan_in_rsci_wen_comp;
  wire [80:0] attenuation_chan_in_rsci_idat_mxwt;
  wire accumalated_color_chan_in_rsci_wen_comp;
  wire [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  wire attenuation_chan_out_rsci_wen_comp;
  reg [80:0] attenuation_chan_out_rsci_idat;
  wire accumalated_color_out_rsci_wen_comp;
  reg [80:0] accumalated_color_out_rsci_idat;
  wire ray_out_loopone_rsci_wen_comp;
  wire ray_out_looptwo_rsci_wen_comp;
  wire ray_out_worldhit_rsci_wen_comp;
  wire quad_out_loopone_rsci_wen_comp;
  reg [376:0] quad_out_loopone_rsci_idat;
  wire quad_out_looptwo_rsci_wen_comp;
  reg [376:0] quad_out_looptwo_rsci_idat;
  wire quad_max_outone_rsci_wen_comp;
  wire quad_max_outtwo_rsci_wen_comp;
  reg [10:0] quad_max_outtwo_rsci_idat;
  wire params_out_rsci_wen_comp;
  reg [92:0] params_out_rsci_idat;
  reg [9:0] quad_max_outone_rsci_idat_9_0;
  wire [9:0] fsm_output;
  wire and_dcpl_2;
  wire and_dcpl_5;
  wire or_tmp_10;
  reg [9:0] reg_params_in_crt_ftd_82;
  reg reg_params_out_rsci_ivld_run_psct_cse;
  wire quad_max_outone_and_cse;
  reg reg_quad_max_outtwo_rsci_ivld_run_psct_cse;
  reg reg_quad_out_looptwo_rsci_ivld_run_psct_cse;
  reg reg_quad_out_loopone_rsci_ivld_run_psct_cse;
  reg reg_ray_out_worldhit_rsci_ivld_run_psct_cse;
  reg [165:0] reg_ray_out_worldhit_rsci_idat_cse;
  reg reg_accumalated_color_out_rsci_ivld_run_psct_cse;
  reg reg_attenuation_chan_out_rsci_ivld_run_psct_cse;
  reg reg_quads_rsci_irdy_run_psct_cse;
  reg reg_params_in_rsci_irdy_run_psct_cse;
  wire params_out_and_cse;
  wire [5:0] for_i_5_0_sva_2;
  wire [6:0] nl_for_i_5_0_sva_2;
  reg for_stage_0_1;
  reg for_stage_0;
  reg [10:0] quad_max_two_sva;
  wire [12:0] nl_quad_max_two_sva;
  reg [4:0] for_i_5_0_sva_4_0;
  wire [10:0] operator_11_false_acc_sdt_sva_1;
  wire [11:0] nl_operator_11_false_acc_sdt_sva_1;

  wire[0:0] or_43_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_LoopDistrib_run_quad_max_outone_rsci_inst_quad_max_outone_rsci_idat;
  assign nl_LoopDistrib_run_quad_max_outone_rsci_inst_quad_max_outone_rsci_idat =
      {1'b0, quad_max_outone_rsci_idat_9_0};
  LoopDistrib_run_ray_in_rsci LoopDistrib_run_ray_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .run_wen(run_wen),
      .ray_in_rsci_oswt(reg_params_out_rsci_ivld_run_psct_cse),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt)
    );
  LoopDistrib_run_params_in_rsci LoopDistrib_run_params_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .run_wen(run_wen),
      .params_in_rsci_oswt(reg_params_in_rsci_irdy_run_psct_cse),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt)
    );
  LoopDistrib_run_quads_rsci LoopDistrib_run_quads_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsc_dat(quads_rsc_dat),
      .quads_rsc_vld(quads_rsc_vld),
      .quads_rsc_rdy(quads_rsc_rdy),
      .run_wen(run_wen),
      .quads_rsci_oswt(reg_quads_rsci_irdy_run_psct_cse),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .quads_rsci_idat_mxwt(quads_rsci_idat_mxwt)
    );
  LoopDistrib_run_attenuation_chan_in_rsci LoopDistrib_run_attenuation_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .run_wen(run_wen),
      .attenuation_chan_in_rsci_oswt(reg_attenuation_chan_out_rsci_ivld_run_psct_cse),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt)
    );
  LoopDistrib_run_accumalated_color_chan_in_rsci LoopDistrib_run_accumalated_color_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .run_wen(run_wen),
      .accumalated_color_chan_in_rsci_oswt(reg_ray_out_worldhit_rsci_ivld_run_psct_cse),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt)
    );
  LoopDistrib_run_attenuation_chan_out_rsci LoopDistrib_run_attenuation_chan_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .run_wen(run_wen),
      .attenuation_chan_out_rsci_oswt(reg_attenuation_chan_out_rsci_ivld_run_psct_cse),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_idat(attenuation_chan_out_rsci_idat)
    );
  LoopDistrib_run_accumalated_color_out_rsci LoopDistrib_run_accumalated_color_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .run_wen(run_wen),
      .accumalated_color_out_rsci_oswt(reg_accumalated_color_out_rsci_ivld_run_psct_cse),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_idat(accumalated_color_out_rsci_idat)
    );
  LoopDistrib_run_ray_out_loopone_rsci LoopDistrib_run_ray_out_loopone_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_loopone_rsc_dat(ray_out_loopone_rsc_dat),
      .ray_out_loopone_rsc_vld(ray_out_loopone_rsc_vld),
      .ray_out_loopone_rsc_rdy(ray_out_loopone_rsc_rdy),
      .run_wen(run_wen),
      .ray_out_loopone_rsci_oswt(reg_ray_out_worldhit_rsci_ivld_run_psct_cse),
      .ray_out_loopone_rsci_wen_comp(ray_out_loopone_rsci_wen_comp),
      .ray_out_loopone_rsci_idat(reg_ray_out_worldhit_rsci_idat_cse)
    );
  LoopDistrib_run_ray_out_looptwo_rsci LoopDistrib_run_ray_out_looptwo_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_looptwo_rsc_dat(ray_out_looptwo_rsc_dat),
      .ray_out_looptwo_rsc_vld(ray_out_looptwo_rsc_vld),
      .ray_out_looptwo_rsc_rdy(ray_out_looptwo_rsc_rdy),
      .run_wen(run_wen),
      .ray_out_looptwo_rsci_oswt(reg_ray_out_worldhit_rsci_ivld_run_psct_cse),
      .ray_out_looptwo_rsci_wen_comp(ray_out_looptwo_rsci_wen_comp),
      .ray_out_looptwo_rsci_idat(reg_ray_out_worldhit_rsci_idat_cse)
    );
  LoopDistrib_run_ray_out_worldhit_rsci LoopDistrib_run_ray_out_worldhit_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_worldhit_rsc_dat(ray_out_worldhit_rsc_dat),
      .ray_out_worldhit_rsc_vld(ray_out_worldhit_rsc_vld),
      .ray_out_worldhit_rsc_rdy(ray_out_worldhit_rsc_rdy),
      .run_wen(run_wen),
      .ray_out_worldhit_rsci_oswt(reg_ray_out_worldhit_rsci_ivld_run_psct_cse),
      .ray_out_worldhit_rsci_wen_comp(ray_out_worldhit_rsci_wen_comp),
      .ray_out_worldhit_rsci_idat(reg_ray_out_worldhit_rsci_idat_cse)
    );
  LoopDistrib_run_quad_out_loopone_rsci LoopDistrib_run_quad_out_loopone_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_out_loopone_rsc_dat(quad_out_loopone_rsc_dat),
      .quad_out_loopone_rsc_vld(quad_out_loopone_rsc_vld),
      .quad_out_loopone_rsc_rdy(quad_out_loopone_rsc_rdy),
      .run_wen(run_wen),
      .quad_out_loopone_rsci_oswt(reg_quad_out_loopone_rsci_ivld_run_psct_cse),
      .quad_out_loopone_rsci_wen_comp(quad_out_loopone_rsci_wen_comp),
      .quad_out_loopone_rsci_idat(quad_out_loopone_rsci_idat)
    );
  LoopDistrib_run_quad_out_looptwo_rsci LoopDistrib_run_quad_out_looptwo_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_out_looptwo_rsc_dat(quad_out_looptwo_rsc_dat),
      .quad_out_looptwo_rsc_vld(quad_out_looptwo_rsc_vld),
      .quad_out_looptwo_rsc_rdy(quad_out_looptwo_rsc_rdy),
      .run_wen(run_wen),
      .quad_out_looptwo_rsci_oswt(reg_quad_out_looptwo_rsci_ivld_run_psct_cse),
      .quad_out_looptwo_rsci_wen_comp(quad_out_looptwo_rsci_wen_comp),
      .quad_out_looptwo_rsci_idat(quad_out_looptwo_rsci_idat)
    );
  LoopDistrib_run_quad_max_outone_rsci LoopDistrib_run_quad_max_outone_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_outone_rsc_dat(quad_max_outone_rsc_dat),
      .quad_max_outone_rsc_vld(quad_max_outone_rsc_vld),
      .quad_max_outone_rsc_rdy(quad_max_outone_rsc_rdy),
      .run_wen(run_wen),
      .quad_max_outone_rsci_oswt(reg_quad_max_outtwo_rsci_ivld_run_psct_cse),
      .quad_max_outone_rsci_wen_comp(quad_max_outone_rsci_wen_comp),
      .quad_max_outone_rsci_idat(nl_LoopDistrib_run_quad_max_outone_rsci_inst_quad_max_outone_rsci_idat[10:0])
    );
  LoopDistrib_run_quad_max_outtwo_rsci LoopDistrib_run_quad_max_outtwo_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_outtwo_rsc_dat(quad_max_outtwo_rsc_dat),
      .quad_max_outtwo_rsc_vld(quad_max_outtwo_rsc_vld),
      .quad_max_outtwo_rsc_rdy(quad_max_outtwo_rsc_rdy),
      .run_wen(run_wen),
      .quad_max_outtwo_rsci_oswt(reg_quad_max_outtwo_rsci_ivld_run_psct_cse),
      .quad_max_outtwo_rsci_wen_comp(quad_max_outtwo_rsci_wen_comp),
      .quad_max_outtwo_rsci_idat(quad_max_outtwo_rsci_idat)
    );
  LoopDistrib_run_params_out_rsci LoopDistrib_run_params_out_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .params_out_rsc_dat(params_out_rsc_dat),
      .params_out_rsc_vld(params_out_rsc_vld),
      .params_out_rsc_rdy(params_out_rsc_rdy),
      .run_wen(run_wen),
      .params_out_rsci_oswt(reg_params_out_rsci_ivld_run_psct_cse),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp),
      .params_out_rsci_idat(params_out_rsci_idat)
    );
  LoopDistrib_run_staller LoopDistrib_run_staller_inst (
      .run_wen(run_wen),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .ray_out_loopone_rsci_wen_comp(ray_out_loopone_rsci_wen_comp),
      .ray_out_looptwo_rsci_wen_comp(ray_out_looptwo_rsci_wen_comp),
      .ray_out_worldhit_rsci_wen_comp(ray_out_worldhit_rsci_wen_comp),
      .quad_out_loopone_rsci_wen_comp(quad_out_loopone_rsci_wen_comp),
      .quad_out_looptwo_rsci_wen_comp(quad_out_looptwo_rsci_wen_comp),
      .quad_max_outone_rsci_wen_comp(quad_max_outone_rsci_wen_comp),
      .quad_max_outtwo_rsci_wen_comp(quad_max_outtwo_rsci_wen_comp),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp)
    );
  LoopDistrib_run_run_fsm LoopDistrib_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_1_tr0(and_dcpl_2)
    );
  assign quad_max_outone_and_cse = run_wen & (~(for_stage_0_1 | for_stage_0 | (~
      (fsm_output[7]))));
  assign params_out_and_cse = run_wen & (fsm_output[1]);
  assign nl_for_i_5_0_sva_2 = conv_u2s_5_6(for_i_5_0_sva_4_0) + 6'b000001;
  assign for_i_5_0_sva_2 = nl_for_i_5_0_sva_2[5:0];
  assign nl_operator_11_false_acc_sdt_sva_1 = conv_u2s_10_11(reg_params_in_crt_ftd_82)
      + 11'b11111111111;
  assign operator_11_false_acc_sdt_sva_1 = nl_operator_11_false_acc_sdt_sva_1[10:0];
  assign and_dcpl_2 = ~(for_stage_0_1 | for_stage_0);
  assign and_dcpl_5 = ~((fsm_output[9]) | (fsm_output[0]));
  assign or_tmp_10 = for_stage_0_1 & (fsm_output[6]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_outone_rsci_idat_9_0 <= 10'b0000000000;
      quad_max_outtwo_rsci_idat <= 11'b00000000000;
    end
    else if ( quad_max_outone_and_cse ) begin
      quad_max_outone_rsci_idat_9_0 <= reg_params_in_crt_ftd_82;
      quad_max_outtwo_rsci_idat <= quad_max_two_sva;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_out_rsci_idat <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quad_max_two_sva <= 11'b00000000000;
    end
    else if ( params_out_and_cse ) begin
      params_out_rsci_idat <= params_in_rsci_idat_mxwt;
      quad_max_two_sva <= nl_quad_max_two_sva[10:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_params_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_quad_max_outtwo_rsci_ivld_run_psct_cse <= 1'b0;
      reg_quad_out_looptwo_rsci_ivld_run_psct_cse <= 1'b0;
      reg_quad_out_loopone_rsci_ivld_run_psct_cse <= 1'b0;
      reg_ray_out_worldhit_rsci_ivld_run_psct_cse <= 1'b0;
      reg_accumalated_color_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_attenuation_chan_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_quads_rsci_irdy_run_psct_cse <= 1'b0;
      reg_params_in_rsci_irdy_run_psct_cse <= 1'b0;
      for_stage_0 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_params_out_rsci_ivld_run_psct_cse <= fsm_output[1];
      reg_quad_max_outtwo_rsci_ivld_run_psct_cse <= and_dcpl_2 & (fsm_output[7]);
      reg_quad_out_looptwo_rsci_ivld_run_psct_cse <= (for_stage_0_1 & (fsm_output[7]))
          | ((quad_max_two_sva[0]) & (fsm_output[8]));
      reg_quad_out_loopone_rsci_ivld_run_psct_cse <= or_tmp_10;
      reg_ray_out_worldhit_rsci_ivld_run_psct_cse <= fsm_output[2];
      reg_accumalated_color_out_rsci_ivld_run_psct_cse <= fsm_output[4];
      reg_attenuation_chan_out_rsci_ivld_run_psct_cse <= fsm_output[3];
      reg_quads_rsci_irdy_run_psct_cse <= ((((~ for_stage_0_1) & (quad_max_two_sva[0]))
          | for_stage_0) & (fsm_output[7])) | (fsm_output[5]) | or_tmp_10;
      reg_params_in_rsci_irdy_run_psct_cse <= ~ and_dcpl_5;
      for_stage_0 <= (for_stage_0 & (~((~((fsm_output[7:6]!=2'b00))) | (((((for_i_5_0_sva_4_0)
          == (operator_11_false_acc_sdt_sva_1[4:0])) & (operator_11_false_acc_sdt_sva_1[10:5]==6'b000000))
          | (for_i_5_0_sva_2[5])) & for_stage_0_1 & (fsm_output[6]))))) | (fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_out_looptwo_rsci_idat <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (~(((~ for_stage_0_1) & (fsm_output[7])) | (~((fsm_output[8:7]!=2'b00)))
        | ((~ (quad_max_two_sva[0])) & (fsm_output[8])))) ) begin
      quad_out_looptwo_rsci_idat <= quads_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_out_loopone_rsci_idat <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[6]) & for_stage_0_1 ) begin
      quad_out_loopone_rsci_idat <= quads_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ray_out_worldhit_rsci_idat_cse <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[2]) ) begin
      reg_ray_out_worldhit_rsci_idat_cse <= ray_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_idat <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[4]) ) begin
      accumalated_color_out_rsci_idat <= attenuation_chan_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_out_rsci_idat <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & (fsm_output[3]) ) begin
      attenuation_chan_out_rsci_idat <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_params_in_crt_ftd_82 <= 10'b0000000000;
    end
    else if ( run_wen & (~(and_dcpl_5 & (~ (fsm_output[1])) & (~ (fsm_output[8]))))
        ) begin
      reg_params_in_crt_ftd_82 <= params_in_rsci_idat_mxwt[10:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_i_5_0_sva_4_0 <= 5'b00000;
    end
    else if ( (for_stage_0_1 | (~ (fsm_output[6]))) & (~ (fsm_output[7])) & run_wen
        ) begin
      for_i_5_0_sva_4_0 <= MUX_v_5_2_2(5'b00000, (for_i_5_0_sva_2[4:0]), (or_43_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_stage_0_1 <= 1'b0;
    end
    else if ( run_wen & ((fsm_output[5]) | (fsm_output[7])) ) begin
      for_stage_0_1 <= for_stage_0 | (fsm_output[5]);
    end
  end
  assign nl_quad_max_two_sva  = (params_in_rsci_idat_mxwt[10:0]) + ({1'b1 , (~ (params_in_rsci_idat_mxwt[10:1]))})
      + 11'b00000000001;
  assign or_43_nl = (fsm_output[7:6]!=2'b00);

  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] conv_u2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_6 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop_hit
// ------------------------------------------------------------------


module IntersecLoop_hit (
  clk, arst_n, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy, ray_temp_in_rsc_dat,
      ray_temp_in_rsc_vld, ray_temp_in_rsc_rdy, quad_max_in_rsc_dat, quad_max_in_rsc_vld,
      quad_max_in_rsc_rdy, quad_hit_anything_out_rsc_dat, quad_hit_anything_out_rsc_vld,
      quad_hit_anything_out_rsc_rdy, rec_quad_out_rsc_dat, rec_quad_out_rsc_vld,
      rec_quad_out_rsc_rdy, closest_so_far_out_rsc_dat, closest_so_far_out_rsc_vld,
      closest_so_far_out_rsc_rdy, mult_run_mul_cmp_a, mult_run_mul_cmp_b, mult_run_mul_cmp_en,
      mult_run_mul_cmp_z, quadInters_qnorm_rorig_run_mul_1_cmp_a, quadInters_qnorm_rorig_run_mul_1_cmp_b,
      quadInters_qnorm_rorig_run_mul_1_cmp_z, quadInters_qnorm_rorig_run_mul_1_cmp_1_a,
      quadInters_qnorm_rorig_run_mul_1_cmp_1_b, quadInters_qnorm_rorig_run_mul_1_cmp_1_z,
      quadInters_qnorm_rorig_run_mul_1_cmp_2_a, quadInters_qnorm_rorig_run_mul_1_cmp_2_b,
      quadInters_qnorm_rorig_run_mul_1_cmp_2_z, quadInters_qnorm_rorig_run_mul_1_cmp_3_a,
      quadInters_qnorm_rorig_run_mul_1_cmp_3_b, quadInters_qnorm_rorig_run_mul_1_cmp_3_z,
      quadInters_qnorm_rorig_run_mul_1_cmp_4_a, quadInters_qnorm_rorig_run_mul_1_cmp_4_b,
      quadInters_qnorm_rorig_run_mul_1_cmp_4_z, quadInters_qnorm_rorig_run_mul_1_cmp_5_a,
      quadInters_qnorm_rorig_run_mul_1_cmp_5_b, quadInters_qnorm_rorig_run_mul_1_cmp_5_z,
      quadInters_denom_dot_run_mul_2_cmp_a, quadInters_denom_dot_run_mul_2_cmp_b,
      quadInters_denom_dot_run_mul_2_cmp_z, quadInters_denom_dot_run_mul_2_cmp_1_a,
      quadInters_denom_dot_run_mul_2_cmp_1_b, quadInters_denom_dot_run_mul_2_cmp_1_z,
      quadInters_denom_dot_run_mul_1_cmp_a, quadInters_denom_dot_run_mul_1_cmp_b,
      quadInters_denom_dot_run_mul_1_cmp_z
);
  input clk;
  input arst_n;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input [165:0] ray_temp_in_rsc_dat;
  input ray_temp_in_rsc_vld;
  output ray_temp_in_rsc_rdy;
  input [10:0] quad_max_in_rsc_dat;
  input quad_max_in_rsc_vld;
  output quad_max_in_rsc_rdy;
  output quad_hit_anything_out_rsc_dat;
  output quad_hit_anything_out_rsc_vld;
  input quad_hit_anything_out_rsc_rdy;
  output [225:0] rec_quad_out_rsc_dat;
  output rec_quad_out_rsc_vld;
  input rec_quad_out_rsc_rdy;
  output [46:0] closest_so_far_out_rsc_dat;
  output closest_so_far_out_rsc_vld;
  input closest_so_far_out_rsc_rdy;
  output [33:0] mult_run_mul_cmp_a;
  output [46:0] mult_run_mul_cmp_b;
  output mult_run_mul_cmp_en;
  input [74:0] mult_run_mul_cmp_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_z;
  output [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_a;
  reg [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_a;
  output [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_b;
  reg [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_b;
  input [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_z;
  output [25:0] quadInters_denom_dot_run_mul_2_cmp_a;
  reg [25:0] quadInters_denom_dot_run_mul_2_cmp_a;
  output [33:0] quadInters_denom_dot_run_mul_2_cmp_b;
  reg [33:0] quadInters_denom_dot_run_mul_2_cmp_b;
  input [57:0] quadInters_denom_dot_run_mul_2_cmp_z;
  output [25:0] quadInters_denom_dot_run_mul_2_cmp_1_a;
  reg [25:0] quadInters_denom_dot_run_mul_2_cmp_1_a;
  output [33:0] quadInters_denom_dot_run_mul_2_cmp_1_b;
  reg [33:0] quadInters_denom_dot_run_mul_2_cmp_1_b;
  input [57:0] quadInters_denom_dot_run_mul_2_cmp_1_z;
  output [25:0] quadInters_denom_dot_run_mul_1_cmp_a;
  reg [25:0] quadInters_denom_dot_run_mul_1_cmp_a;
  output [33:0] quadInters_denom_dot_run_mul_1_cmp_b;
  reg [33:0] quadInters_denom_dot_run_mul_1_cmp_b;
  input [59:0] quadInters_denom_dot_run_mul_1_cmp_z;


  // Interconnect Declarations
  wire hit_wen;
  wire quads_rsci_wen_comp;
  wire [376:0] quads_rsci_idat_mxwt;
  wire ray_temp_in_rsci_wen_comp;
  wire [165:0] ray_temp_in_rsci_idat_mxwt;
  wire quad_max_in_rsci_wen_comp;
  wire [10:0] quad_max_in_rsci_idat_mxwt;
  wire quad_hit_anything_out_rsci_wen_comp;
  reg quad_hit_anything_out_rsci_idat;
  wire rec_quad_out_rsci_wen_comp;
  wire closest_so_far_out_rsci_wen_comp;
  reg ensig_cgo;
  wire [44:0] mult_run_mul_cmp_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg;
  wire [61:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg;
  wire [57:0] quadInters_denom_dot_run_mul_2_cmp_z_oreg;
  wire [57:0] quadInters_denom_dot_run_mul_2_cmp_1_z_oreg;
  wire [59:0] quadInters_denom_dot_run_mul_1_cmp_z_oreg;
  reg [26:0] rec_quad_out_rsci_idat_225_199;
  reg [26:0] rec_quad_out_rsci_idat_198_172;
  reg [26:0] rec_quad_out_rsci_idat_171_145;
  reg [2:0] rec_quad_out_rsci_idat_144_142;
  reg rec_quad_out_rsci_idat_141;
  reg [25:0] rec_quad_out_rsci_idat_140_115;
  reg [25:0] rec_quad_out_rsci_idat_114_89;
  reg [25:0] rec_quad_out_rsci_idat_88_63;
  reg [19:0] rec_quad_out_rsci_idat_62_43;
  reg rec_quad_out_rsci_idat_42;
  reg [19:0] rec_quad_out_rsci_idat_41_22;
  reg rec_quad_out_rsci_idat_21;
  reg [19:0] rec_quad_out_rsci_idat_20_1;
  reg rec_quad_out_rsci_idat_0;
  reg closest_so_far_out_rsci_idat_46;
  reg closest_so_far_out_rsci_idat_45;
  reg closest_so_far_out_rsci_idat_44;
  reg closest_so_far_out_rsci_idat_43;
  reg closest_so_far_out_rsci_idat_42;
  reg closest_so_far_out_rsci_idat_41;
  reg closest_so_far_out_rsci_idat_40;
  reg closest_so_far_out_rsci_idat_39;
  reg closest_so_far_out_rsci_idat_38;
  reg closest_so_far_out_rsci_idat_37;
  reg closest_so_far_out_rsci_idat_36;
  reg closest_so_far_out_rsci_idat_35;
  reg closest_so_far_out_rsci_idat_34;
  reg closest_so_far_out_rsci_idat_33;
  reg closest_so_far_out_rsci_idat_32;
  reg closest_so_far_out_rsci_idat_31;
  reg closest_so_far_out_rsci_idat_30;
  reg closest_so_far_out_rsci_idat_29;
  reg closest_so_far_out_rsci_idat_28;
  reg closest_so_far_out_rsci_idat_27;
  reg closest_so_far_out_rsci_idat_26;
  reg closest_so_far_out_rsci_idat_25;
  reg closest_so_far_out_rsci_idat_24;
  reg closest_so_far_out_rsci_idat_23;
  reg closest_so_far_out_rsci_idat_22;
  reg closest_so_far_out_rsci_idat_21;
  reg closest_so_far_out_rsci_idat_20;
  reg closest_so_far_out_rsci_idat_19;
  reg closest_so_far_out_rsci_idat_18;
  reg closest_so_far_out_rsci_idat_17;
  reg closest_so_far_out_rsci_idat_16;
  reg closest_so_far_out_rsci_idat_15;
  reg closest_so_far_out_rsci_idat_14;
  reg closest_so_far_out_rsci_idat_13;
  reg closest_so_far_out_rsci_idat_12;
  reg closest_so_far_out_rsci_idat_11;
  reg closest_so_far_out_rsci_idat_10;
  reg closest_so_far_out_rsci_idat_9;
  reg closest_so_far_out_rsci_idat_8;
  reg closest_so_far_out_rsci_idat_7;
  reg closest_so_far_out_rsci_idat_6;
  reg closest_so_far_out_rsci_idat_5;
  reg closest_so_far_out_rsci_idat_4;
  reg closest_so_far_out_rsci_idat_3;
  reg closest_so_far_out_rsci_idat_2;
  reg closest_so_far_out_rsci_idat_1;
  reg closest_so_far_out_rsci_idat_0;
  wire [6:0] fsm_output;
  wire for_nor_tmp;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp;
  wire quadInters_run_if_5_quadInters_run_if_5_or_2_tmp;
  wire and_dcpl_54;
  wire and_dcpl_195;
  wire or_dcpl_79;
  wire and_dcpl_200;
  wire or_dcpl_91;
  wire or_dcpl_95;
  wire and_dcpl_238;
  wire or_tmp_328;
  wire or_tmp_480;
  wire or_tmp_481;
  wire or_tmp_490;
  wire or_tmp_529;
  wire or_tmp_531;
  wire or_tmp_673;
  wire or_tmp_691;
  wire quadInters_run_mux_593_tmp_33;
  wire and_1128_cse;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_33_itm;
  reg quadInters_run_lor_3_lpi_2_dfm_1;
  reg quadInters_run_lor_lpi_2_dfm_2;
  wire quadInters_run_or_1_tmp_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm;
  reg quadInters_run_land_lpi_2_dfm_9;
  reg quadInters_run_lor_lpi_2_dfm_1;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7;
  reg quadInters_run_land_lpi_2_dfm_8;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_2_itm_1;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm;
  reg quadInters_run_lor_lpi_2_dfm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_33_itm;
  reg for_stage_0_9;
  reg for_hitWorld_lpi_2_dfm_2;
  reg for_stage_0_3;
  reg quadInters_run_land_lpi_2_dfm_st_2;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_1;
  reg for_stage_0_4;
  reg quadInters_run_land_lpi_2_dfm_st_3;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2;
  reg for_stage_0_5;
  reg quadInters_run_land_lpi_2_dfm_st_4;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3;
  reg for_stage_0_6;
  reg quadInters_run_land_lpi_2_dfm_st_5;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_4;
  reg for_stage_0_7;
  reg quadInters_run_land_lpi_2_dfm_st_6;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_5;
  reg quadInters_run_lor_3_lpi_2_dfm;
  reg [165:0] ray_temp_in_crt_sva;
  reg for_stage_0_2;
  reg quadInters_run_land_lpi_2_dfm_st_1;
  reg for_stage_0_8;
  reg quadInters_run_land_lpi_2_dfm_st_7;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_1_itm;
  reg for_stage_0_1;
  reg for_stage_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4;
  reg quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st;
  reg operator_33_true_asn_1_itm_9;
  reg operator_33_true_asn_1_itm_7;
  reg operator_33_true_asn_1_itm_8;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_1;
  reg quadInters_run_land_lpi_2_dfm;
  reg [59:0] setfacenorm_dot_run_acc_2_itm;
  reg [4:0] for_i_5_0_sva_4_0;
  wire [11:0] operator_11_false_acc_sdt_sva_1;
  wire [12:0] nl_operator_11_false_acc_sdt_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_73_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_74_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_68_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_mx2;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_50_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_40_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx3;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1;
  wire [1:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx0_33_32;
  wire ensig_cgo_mx0;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd;
  reg [32:0] reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd_1;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd;
  reg [32:0] reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd;
  reg reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1;
  wire closest_so_far_out_and_cse;
  reg reg_closest_so_far_out_rsci_ivld_hit_psct_cse;
  reg reg_quad_max_in_rsci_irdy_hit_psct_cse;
  reg reg_quads_rsci_irdy_hit_psct_cse;
  wire closest_so_far_and_cse;
  wire or_343_cse;
  wire for_and_1_cse;
  wire or_69_cse;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_46;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_45;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_44;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_43;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_42;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_41;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_40;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_39;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_38;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_37;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_36;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_35;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_34;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_33;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_32;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_31;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_30;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_29;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_28;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_27;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_26;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_25;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_24;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_23;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_22;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_21;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_20;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_19;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_18;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_17;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_16;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_15;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_14;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_13;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_12;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_11;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_10;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_9;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_8;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_7;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_6;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_5;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_4;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_3;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_2;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_1;
  reg quadInters_run_t_trunc_lpi_2_dfm_1_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  wire quadInters_run_t_trunc_lpi_2_dfm_45_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_44_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_43_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_42_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_41_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_40_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_39_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_38_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_37_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_36_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_35_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_34_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_33_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_32_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_31_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_30_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_29_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_28_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_27_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_26_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_25_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_24_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_23_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_22_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_21_1;
  wire quadInters_run_t_trunc_lpi_2_dfm_20_1;
  wire and_454_cse;
  reg [80:0] quads_crt_sva_8_376_296;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_mux_10_itm;
  wire [59:0] z_out;
  wire [20:0] z_out_1;
  wire [21:0] nl_z_out_1;
  wire [33:0] z_out_2;
  wire [34:0] nl_z_out_2;
  wire [34:0] z_out_3;
  wire [35:0] nl_z_out_3;
  wire [33:0] z_out_4;
  wire [34:0] nl_z_out_4;
  wire [33:0] z_out_5;
  wire [34:0] nl_z_out_5;
  wire [33:0] z_out_6;
  wire [34:0] nl_z_out_6;
  wire [33:0] z_out_7;
  wire [34:0] nl_z_out_7;
  wire [34:0] z_out_8;
  wire [35:0] nl_z_out_8;
  wire [34:0] z_out_9;
  wire [35:0] nl_z_out_9;
  wire [34:0] z_out_10;
  wire [35:0] nl_z_out_10;
  wire [34:0] z_out_11;
  wire [35:0] nl_z_out_11;
  wire [34:0] z_out_12;
  wire [35:0] nl_z_out_12;
  wire [34:0] z_out_13;
  wire [35:0] nl_z_out_13;
  wire [34:0] z_out_14;
  wire [35:0] nl_z_out_14;
  reg [25:0] quadInters_setfacenorm_run_qr_x_lpi_2;
  reg [25:0] quadInters_setfacenorm_run_qr_y_lpi_2;
  reg [25:0] quadInters_setfacenorm_run_qr_z_lpi_2;
  reg [10:0] quad_max_sva;
  reg quad_hit_anything_sva;
  reg rec_quad_hit_loc_x_0_sva;
  reg [19:0] rec_quad_hit_loc_x_20_1_sva;
  reg rec_quad_hit_loc_y_0_sva;
  reg [19:0] rec_quad_hit_loc_y_20_1_sva;
  reg rec_quad_hit_loc_z_0_sva;
  reg [19:0] rec_quad_hit_loc_z_20_1_sva;
  reg [25:0] rec_quad_normal_x_sva;
  reg [25:0] rec_quad_normal_y_sva;
  reg [25:0] rec_quad_normal_z_sva;
  reg rec_quad_front_face_sva;
  reg [2:0] rec_quad_mat_sva;
  reg [26:0] rec_quad_color_r_sva;
  reg [26:0] rec_quad_color_g_sva;
  reg [26:0] rec_quad_color_b_sva;
  reg [376:0] quads_crt_sva;
  reg [33:0] ac_math_ac_abs_58_58_xabs_57_24_sva;
  reg [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva;
  reg [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_57_lpi_2_dfm;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm;
  reg [31:0] add_run_ac_fixed_cctor_74_43_sva;
  reg [31:0] add_run_ac_fixed_cctor_1_74_43_sva;
  reg [31:0] add_run_ac_fixed_cctor_2_74_43_sva;
  reg quad_hit_anything_sva_dfm;
  reg [25:0] rec_quad_normal_x_sva_dfm;
  reg [25:0] rec_quad_normal_y_sva_dfm;
  reg [25:0] rec_quad_normal_z_sva_dfm;
  reg [26:0] rec_quad_color_r_sva_dfm;
  reg [26:0] rec_quad_color_g_sva_dfm;
  reg [26:0] rec_quad_color_b_sva_dfm;
  reg rec_quad_hit_loc_x_0_sva_dfm;
  reg rec_quad_hit_loc_y_0_sva_dfm;
  reg rec_quad_hit_loc_z_0_sva_dfm;
  reg [57:0] ac_math_ac_abs_58_58_xabs_xor_itm;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_itm;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_33_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_46_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_47_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_33_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_33_itm;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_33_itm;
  reg operator_33_true_asn_1_itm;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3;
  reg [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_6_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_5_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_4_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_3_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_33_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_33_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_9_psp_33_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_33_itm_1;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1;
  reg operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_33_itm_1;
  reg operator_33_true_asn_1_itm_1;
  reg operator_33_true_asn_1_itm_2;
  reg operator_33_true_asn_1_itm_3;
  reg operator_33_true_asn_1_itm_4;
  reg operator_33_true_asn_1_itm_5;
  reg operator_33_true_asn_1_itm_6;
  reg closest_so_far_sva_46;
  reg closest_so_far_sva_45;
  reg closest_so_far_sva_44;
  reg closest_so_far_sva_43;
  reg closest_so_far_sva_42;
  reg closest_so_far_sva_41;
  reg closest_so_far_sva_40;
  reg closest_so_far_sva_39;
  reg closest_so_far_sva_38;
  reg closest_so_far_sva_37;
  reg closest_so_far_sva_36;
  reg closest_so_far_sva_35;
  reg closest_so_far_sva_34;
  reg closest_so_far_sva_33;
  reg closest_so_far_sva_32;
  reg closest_so_far_sva_31;
  reg closest_so_far_sva_30;
  reg closest_so_far_sva_29;
  reg closest_so_far_sva_28;
  reg closest_so_far_sva_27;
  reg closest_so_far_sva_26;
  reg closest_so_far_sva_25;
  reg closest_so_far_sva_24;
  reg closest_so_far_sva_23;
  reg closest_so_far_sva_22;
  reg closest_so_far_sva_21;
  reg closest_so_far_sva_20;
  reg closest_so_far_sva_19;
  reg closest_so_far_sva_18;
  reg closest_so_far_sva_17;
  reg closest_so_far_sva_16;
  reg closest_so_far_sva_15;
  reg closest_so_far_sva_14;
  reg closest_so_far_sva_13;
  reg closest_so_far_sva_12;
  reg closest_so_far_sva_11;
  reg closest_so_far_sva_10;
  reg closest_so_far_sva_9;
  reg closest_so_far_sva_8;
  reg closest_so_far_sva_7;
  reg closest_so_far_sva_6;
  reg closest_so_far_sva_5;
  reg closest_so_far_sva_4;
  reg closest_so_far_sva_3;
  reg closest_so_far_sva_2;
  reg closest_so_far_sva_1;
  reg closest_so_far_sva_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_45;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_44;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_43;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_42;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_41;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_40;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_39;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_38;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_37;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_36;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_35;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_34;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_32;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_31;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_30;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_29;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_28;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_27;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_26;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_25;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_24;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_23;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_22;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_21;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_9;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_8;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_7;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_6;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_5;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_4;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_3;
  reg closest_so_far_sva_dfm_3_46;
  reg closest_so_far_sva_dfm_3_45;
  reg closest_so_far_sva_dfm_3_44;
  reg closest_so_far_sva_dfm_3_43;
  reg closest_so_far_sva_dfm_3_42;
  reg closest_so_far_sva_dfm_3_41;
  reg closest_so_far_sva_dfm_3_40;
  reg closest_so_far_sva_dfm_3_39;
  reg closest_so_far_sva_dfm_3_38;
  reg closest_so_far_sva_dfm_3_37;
  reg closest_so_far_sva_dfm_3_36;
  reg closest_so_far_sva_dfm_3_35;
  reg closest_so_far_sva_dfm_3_34;
  reg closest_so_far_sva_dfm_3_33;
  reg closest_so_far_sva_dfm_3_32;
  reg closest_so_far_sva_dfm_3_31;
  reg closest_so_far_sva_dfm_3_30;
  reg closest_so_far_sva_dfm_3_29;
  reg closest_so_far_sva_dfm_3_28;
  reg closest_so_far_sva_dfm_3_27;
  reg closest_so_far_sva_dfm_3_26;
  reg closest_so_far_sva_dfm_3_25;
  reg closest_so_far_sva_dfm_3_24;
  reg closest_so_far_sva_dfm_3_23;
  reg closest_so_far_sva_dfm_3_22;
  reg closest_so_far_sva_dfm_3_21;
  reg closest_so_far_sva_dfm_3_20;
  reg closest_so_far_sva_dfm_3_19;
  reg closest_so_far_sva_dfm_3_18;
  reg closest_so_far_sva_dfm_3_17;
  reg closest_so_far_sva_dfm_3_16;
  reg closest_so_far_sva_dfm_3_15;
  reg closest_so_far_sva_dfm_3_14;
  reg closest_so_far_sva_dfm_3_13;
  reg closest_so_far_sva_dfm_3_12;
  reg closest_so_far_sva_dfm_3_11;
  reg closest_so_far_sva_dfm_3_10;
  reg closest_so_far_sva_dfm_3_9;
  reg closest_so_far_sva_dfm_3_8;
  reg closest_so_far_sva_dfm_3_7;
  reg closest_so_far_sva_dfm_3_6;
  reg closest_so_far_sva_dfm_3_5;
  reg closest_so_far_sva_dfm_3_4;
  reg closest_so_far_sva_dfm_3_3;
  reg closest_so_far_sva_dfm_3_2;
  reg closest_so_far_sva_dfm_3_1;
  reg closest_so_far_sva_dfm_3_0;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_46;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_45;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_44;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_43;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_42;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_41;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_40;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_39;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_38;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_37;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_36;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_35;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_34;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_33;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_32;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_31;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_30;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_29;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_28;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_27;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_26;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_25;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_24;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_23;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_22;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_21;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_20;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_19;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_18;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_17;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_16;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_15;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_14;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_13;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_12;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_11;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_10;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_9;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_8;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_7;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_6;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_5;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_4;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_3;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_2;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_1;
  reg quadInters_run_t_trunc_lpi_2_dfm_2_0;
  reg [264:0] quads_crt_sva_1_376_112;
  reg [110:0] quads_crt_sva_1_110_0;
  reg [80:0] quads_crt_sva_2_376_296;
  reg [152:0] quads_crt_sva_2_264_112;
  reg [110:0] quads_crt_sva_2_110_0;
  reg [80:0] quads_crt_sva_3_376_296;
  reg [152:0] quads_crt_sva_3_264_112;
  reg [110:0] quads_crt_sva_3_110_0;
  reg [80:0] quads_crt_sva_4_376_296;
  reg [152:0] quads_crt_sva_4_264_112;
  reg [110:0] quads_crt_sva_4_110_0;
  reg [80:0] quads_crt_sva_5_376_296;
  reg [152:0] quads_crt_sva_5_264_112;
  reg [110:0] quads_crt_sva_5_110_0;
  reg [80:0] quads_crt_sva_6_376_296;
  reg [152:0] quads_crt_sva_6_264_112;
  reg [110:0] quads_crt_sva_6_110_0;
  reg [80:0] quads_crt_sva_7_376_296;
  reg [152:0] quads_crt_sva_7_264_112;
  reg [110:0] quads_crt_sva_7_110_0;
  reg [77:0] quads_crt_sva_8_189_112;
  reg [2:0] quads_crt_sva_8_110_108;
  reg [77:0] quads_crt_sva_9_189_112;
  reg [44:0] mult_run_asn_2_itm_1_74_30;
  wire quad_hit_anything_sva_dfm_mx0w0;
  wire quadInters_run_quadInters_run_quadInters_run_nor_6_mx0w1;
  wire [19:0] quadInters_run_quadInters_run_and_6_mx0w2;
  wire quadInters_run_quadInters_run_quadInters_run_nor_5_mx0w1;
  wire [19:0] quadInters_run_quadInters_run_and_4_mx0w2;
  wire quadInters_run_quadInters_run_quadInters_run_nor_mx0w1;
  wire [19:0] quadInters_run_quadInters_run_and_2_mx0w2;
  wire [31:0] add_run_ac_fixed_cctor_2_74_43_sva_mx1w0;
  wire [32:0] nl_add_run_ac_fixed_cctor_2_74_43_sva_mx1w0;
  wire [31:0] add_run_ac_fixed_cctor_1_74_43_sva_mx1w0;
  wire [32:0] nl_add_run_ac_fixed_cctor_1_74_43_sva_mx1w0;
  wire [31:0] add_run_ac_fixed_cctor_74_43_sva_mx1w0;
  wire [32:0] nl_add_run_ac_fixed_cctor_74_43_sva_mx1w0;
  wire quadInters_run_lor_lpi_2_dfm_mx0w1;
  wire operator_33_true_asn_1_itm_9_mx0c2;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0;
  wire [25:0] quadInters_setfacenorm_run_qr_z_lpi_2_dfm_4_mx1w0;
  wire [25:0] quadInters_setfacenorm_run_qr_y_lpi_2_dfm_4_mx1w0;
  wire [25:0] quadInters_setfacenorm_run_qr_x_lpi_2_dfm_4_mx1w0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx2;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_mx1w0;
  wire for_hitWorld_lpi_2_dfm_3;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_72_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_71_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_70_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_69_lpi_2_dfm_mx0;
  wire [33:0] ac_math_ac_abs_58_58_xabs_57_24_sva_mx1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_49_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_48_lpi_2_dfm_mx0;
  wire [57:0] quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0;
  wire [58:0] nl_quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0;
  wire quadInters_run_quadInters_run_nor_4_cse_1;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_77_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_76_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_75_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_55_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_54_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_53_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_52_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_35_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_34_lpi_2_dfm_mx0;
  wire quadInters_run_asn_69;
  wire quadInters_run_asn_71;
  wire [34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2;
  wire [35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_lpi_2_dfm_34_1_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_60_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_59_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_58_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_39_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_38_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_66_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_65_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_64_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_63_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_46_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_45_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_44_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_43_lpi_2_dfm_mx0;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_42_lpi_2_dfm_mx0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_18_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_20_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_33;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_0;
  reg [12:0] quadInters_at_run_mult_result_x_74_30_sva_12_0;
  wire [32:0] quadInters_run_rounded_denom_lpi_2_dfm_mx0_32_0;
  wire [1:0] quadInters_run_if_1_exs_mx1w0_1_0;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_qelse_conc_itm_33;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_m1c;
  reg [19:0] reg_ac_math_ac_abs_21_21_xabs_xor_ftd_1;
  reg [19:0] reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1;
  reg [19:0] reg_ac_math_ac_abs_21_21_1_xabs_xor_ftd_1;
  wire rec_quad_mat_and_1_rgt;
  wire quadInters_denom_dot_run_and_4_rgt;
  wire quadInters_denom_dot_run_and_5_rgt;
  wire operator_35_true_and_30_rgt;
  wire operator_35_true_and_31_rgt;
  wire operator_35_true_and_32_rgt;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_6_rgt;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_or_rgt;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_rgt;
  wire operator_35_true_and_16_rgt;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_and_rgt;
  wire operator_35_true_and_57_cse;
  wire operator_35_true_and_58_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_12_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_13_cse;
  wire quadInters_run_t_trunc_mux_47_cse;
  wire quadInters_run_t_trunc_mux_48_cse;
  wire quadInters_run_t_trunc_mux_49_cse;
  wire quadInters_run_t_trunc_mux_50_cse;
  wire quadInters_run_t_trunc_mux_51_cse;
  wire quadInters_run_t_trunc_mux_52_cse;
  wire quadInters_run_t_trunc_mux_53_cse;
  wire quadInters_run_t_trunc_mux_54_cse;
  wire quadInters_run_t_trunc_mux_55_cse;
  wire quadInters_run_t_trunc_mux_56_cse;
  wire quadInters_run_t_trunc_mux_57_cse;
  wire quadInters_run_t_trunc_mux_58_cse;
  wire quadInters_run_t_trunc_mux_59_cse;
  wire quadInters_run_t_trunc_mux_60_cse;
  wire quadInters_run_t_trunc_mux_61_cse;
  wire quadInters_run_t_trunc_mux_62_cse;
  wire quadInters_run_t_trunc_mux_63_cse;
  wire quadInters_run_t_trunc_mux_64_cse;
  wire quadInters_run_t_trunc_mux_65_cse;
  wire quadInters_run_t_trunc_mux_66_cse;
  wire quadInters_run_t_trunc_mux_67_cse;
  wire quadInters_run_t_trunc_mux_68_cse;
  wire quadInters_run_t_trunc_mux_69_cse;
  wire quadInters_run_t_trunc_mux_70_cse;
  wire quadInters_run_t_trunc_mux_71_cse;
  wire quadInters_run_t_trunc_mux_72_cse;
  wire quadInters_run_t_trunc_mux_73_cse;
  wire quadInters_run_t_trunc_mux_74_cse;
  wire quadInters_run_t_trunc_mux_75_cse;
  wire quadInters_run_t_trunc_mux_76_cse;
  wire quadInters_run_t_trunc_mux_77_cse;
  wire quadInters_run_t_trunc_mux_78_cse;
  wire quadInters_run_t_trunc_mux_79_cse;
  wire quadInters_run_t_trunc_mux_80_cse;
  wire quadInters_run_t_trunc_mux_81_cse;
  wire quadInters_run_t_trunc_mux_82_cse;
  wire quadInters_run_t_trunc_mux_83_cse;
  wire quadInters_run_t_trunc_mux_84_cse;
  wire quadInters_run_t_trunc_mux_85_cse;
  wire quadInters_run_t_trunc_mux_86_cse;
  wire quadInters_run_t_trunc_mux_87_cse;
  wire quadInters_run_t_trunc_mux_88_cse;
  wire quadInters_run_t_trunc_mux_89_cse;
  wire quadInters_run_t_trunc_mux_90_cse;
  wire quadInters_run_t_trunc_mux_91_cse;
  wire quadInters_run_t_trunc_mux_92_cse;
  wire quadInters_run_t_trunc_mux_93_cse;
  wire closest_so_far_and_47_cse;
  wire rec_quad_color_b_and_cse;
  wire rec_quad_normal_z_and_cse;
  wire rec_quad_hit_loc_z_and_cse;
  wire add_run_and_3_cse;
  wire ac_math_ac_abs_21_21_1_xabs_and_1_cse;
  wire quadInters_run_oelse_and_1_cse;
  wire operator_35_true_and_59_cse;
  wire operator_35_true_and_100_cse;
  wire operator_35_true_and_282_cse;
  wire operator_35_true_and_135_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_cse;
  wire quadInters_run_oelse_and_2_cse;
  wire operator_35_true_and_185_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_1_cse;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_5_cse;
  reg reg_quadInters_run_if_4_slc_quadInters_run_if_4_acc_27_svs_st_1_cse;
  wire [33:0] quadInters_denom_dot_run_mux1h_5_rgt;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_11_rgt;
  wire [22:0] quadInters_sub_run_mux_rgt;
  wire [22:0] quadInters_sub_run_mux_1_rgt;
  wire [22:0] quadInters_sub_run_mux_2_rgt;
  wire [33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt;
  wire [34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33;
  reg [32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_32_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33;
  reg [32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_32_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33;
  reg [1:0] quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56;
  reg [31:0] quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24;
  reg [4:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22;
  reg [21:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0;
  reg [33:0] quadInters_denom_dot_run_ac_fixed_cctor_sva_57_24;
  reg [23:0] quadInters_denom_dot_run_ac_fixed_cctor_sva_23_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33;
  reg [32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_32_0;
  reg div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33;
  reg [32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_32_0;
  reg [31:0] mult_run_asn_1_itm_74_43;
  reg [12:0] mult_run_asn_1_itm_42_30;
  reg [1:0] reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg;
  reg [20:0] reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg;
  reg [1:0] reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg;
  reg [20:0] reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg;
  reg [1:0] reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg;
  reg [20:0] reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg;
  wire and_2744_cse;
  wire and_2754_cse;
  wire and_2778_cse;
  wire and_1706_cse;
  wire and_2843_cse;
  wire and_2862_cse;
  wire and_2865_cse;
  wire or_1462_cse;
  wire or_cse;
  reg [32:0] reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_1_cse;
  wire and_2828_cse;
  wire operator_38_15_true_AC_TRN_AC_WRAP_1_acc_itm_38;
  wire operator_38_15_true_AC_TRN_AC_WRAP_acc_itm_38;
  wire [37:0] quadInters_beta_dot_run_acc_itm_61_24;
  wire [37:0] quadInters_alpha_dot_run_acc_itm_61_24;
  wire [33:0] ac_math_ac_abs_58_58_xabs_acc_itm_57_24;
  wire setfacenorm_dot_run_acc_itm_59;
  wire quadInters_run_acc_6_itm_21;
  wire quadInters_run_acc_5_itm_21;
  wire quadInters_run_acc_4_itm_21;
  wire [46:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13;
  wire quadInters_run_if_1_acc_itm_34;
  wire div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_3_cse;

  wire[56:0] quadInters_cross_u_run_acc_nl;
  wire[57:0] nl_quadInters_cross_u_run_acc_nl;
  wire[56:0] quadInters_cross_u_run_mul_nl;
  wire[56:0] quadInters_cross_u_run_mul_1_nl;
  wire[56:0] quadInters_cross_u_run_acc_2_nl;
  wire[57:0] nl_quadInters_cross_u_run_acc_2_nl;
  wire[56:0] quadInters_cross_u_run_mul_4_nl;
  wire[56:0] quadInters_cross_u_run_mul_5_nl;
  wire[56:0] quadInters_cross_v_run_acc_2_nl;
  wire[57:0] nl_quadInters_cross_v_run_acc_2_nl;
  wire[56:0] quadInters_cross_v_run_mul_4_nl;
  wire[56:0] quadInters_cross_v_run_mul_5_nl;
  wire[56:0] quadInters_cross_v_run_acc_nl;
  wire[57:0] nl_quadInters_cross_v_run_acc_nl;
  wire[56:0] quadInters_cross_v_run_mul_nl;
  wire[56:0] quadInters_cross_v_run_mul_1_nl;
  wire[56:0] quadInters_cross_u_run_acc_1_nl;
  wire[57:0] nl_quadInters_cross_u_run_acc_1_nl;
  wire[56:0] quadInters_cross_u_run_mul_2_nl;
  wire[56:0] quadInters_cross_u_run_mul_3_nl;
  wire[19:0] rec_quad_hit_loc_x_asn_ac_math_ac_abs_21_21_1_xabs_xor_itm_mx1w1_19_and_nl;
  wire[19:0] mux_125_nl;
  wire[0:0] not_nl;
  wire[19:0] ac_math_ac_abs_21_21_1_xabs_xor_1_nl;
  wire[19:0] rec_quad_hit_loc_y_asn_ac_math_ac_abs_21_21_2_xabs_xor_itm_mx1w1_19_and_nl;
  wire[19:0] mux_124_nl;
  wire[0:0] not_669_nl;
  wire[19:0] ac_math_ac_abs_21_21_2_xabs_xor_1_nl;
  wire[19:0] rec_quad_hit_loc_z_asn_ac_math_ac_abs_21_21_xabs_xor_itm_mx1w1_19_and_nl;
  wire[19:0] mux_123_nl;
  wire[0:0] not_670_nl;
  wire[19:0] ac_math_ac_abs_21_21_xabs_xor_1_nl;
  wire[0:0] quad_hit_anything_mux_48_nl;
  wire[0:0] quad_hit_anything_mux_47_nl;
  wire[0:0] quad_hit_anything_mux_46_nl;
  wire[0:0] quad_hit_anything_mux_45_nl;
  wire[0:0] quad_hit_anything_mux_44_nl;
  wire[0:0] quad_hit_anything_mux_43_nl;
  wire[0:0] quad_hit_anything_mux_42_nl;
  wire[0:0] quad_hit_anything_mux_41_nl;
  wire[0:0] quad_hit_anything_mux_40_nl;
  wire[0:0] quad_hit_anything_mux_39_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_4_nl;
  wire[0:0] quad_hit_anything_mux_38_nl;
  wire[0:0] quad_hit_anything_mux_37_nl;
  wire[0:0] quad_hit_anything_mux_36_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_3_nl;
  wire[0:0] quad_hit_anything_mux_35_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_2_nl;
  wire[0:0] quad_hit_anything_mux_34_nl;
  wire[0:0] quad_hit_anything_mux_33_nl;
  wire[0:0] quad_hit_anything_mux_32_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_1_nl;
  wire[0:0] quad_hit_anything_mux_31_nl;
  wire[0:0] quad_hit_anything_mux_30_nl;
  wire[0:0] quad_hit_anything_mux_29_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_nl;
  wire[0:0] quad_hit_anything_mux_28_nl;
  wire[0:0] quad_hit_anything_mux_27_nl;
  wire[0:0] quad_hit_anything_mux_26_nl;
  wire[0:0] quad_hit_anything_mux_25_nl;
  wire[0:0] quad_hit_anything_mux_24_nl;
  wire[0:0] quad_hit_anything_mux_23_nl;
  wire[0:0] quad_hit_anything_mux_22_nl;
  wire[0:0] quad_hit_anything_mux_21_nl;
  wire[0:0] quad_hit_anything_mux_20_nl;
  wire[0:0] quad_hit_anything_mux_19_nl;
  wire[0:0] quad_hit_anything_mux_18_nl;
  wire[0:0] quad_hit_anything_mux_17_nl;
  wire[0:0] quad_hit_anything_mux_16_nl;
  wire[0:0] quad_hit_anything_mux_15_nl;
  wire[0:0] quad_hit_anything_mux_14_nl;
  wire[0:0] quad_hit_anything_mux_13_nl;
  wire[0:0] quad_hit_anything_mux_12_nl;
  wire[0:0] quad_hit_anything_mux_11_nl;
  wire[0:0] quad_hit_anything_mux_10_nl;
  wire[0:0] quad_hit_anything_mux_9_nl;
  wire[0:0] quad_hit_anything_mux_8_nl;
  wire[0:0] quad_hit_anything_mux_7_nl;
  wire[0:0] quad_hit_anything_mux_6_nl;
  wire[0:0] not_676_nl;
  wire[0:0] quad_hit_anything_mux_5_nl;
  wire[0:0] not_674_nl;
  wire[0:0] quad_hit_anything_mux_4_nl;
  wire[0:0] not_672_nl;
  wire[0:0] rec_quad_color_b_not_nl;
  wire[0:0] rec_quad_color_g_not_nl;
  wire[0:0] rec_quad_color_r_not_nl;
  wire[0:0] rec_quad_mat_not_nl;
  wire[0:0] quad_hit_anything_mux_nl;
  wire[0:0] quad_hit_anything_mux_2_nl;
  wire[0:0] quadInters_run_quadInters_run_or_10_nl;
  wire[0:0] quadInters_run_quadInters_run_or_12_nl;
  wire[0:0] quadInters_run_quadInters_run_or_14_nl;
  wire[0:0] quadInters_run_quadInters_run_or_16_nl;
  wire[0:0] quadInters_run_quadInters_run_or_18_nl;
  wire[0:0] quadInters_run_quadInters_run_or_20_nl;
  wire[0:0] quadInters_run_quadInters_run_or_22_nl;
  wire[0:0] quadInters_run_quadInters_run_or_24_nl;
  wire[0:0] quadInters_run_quadInters_run_or_26_nl;
  wire[0:0] quadInters_run_quadInters_run_or_28_nl;
  wire[0:0] quadInters_run_quadInters_run_or_30_nl;
  wire[0:0] quadInters_run_quadInters_run_or_32_nl;
  wire[0:0] quadInters_run_quadInters_run_or_34_nl;
  wire[0:0] quadInters_run_quadInters_run_or_36_nl;
  wire[0:0] quadInters_run_quadInters_run_or_38_nl;
  wire[0:0] quadInters_run_quadInters_run_or_40_nl;
  wire[0:0] quadInters_run_quadInters_run_or_42_nl;
  wire[0:0] quadInters_run_quadInters_run_or_44_nl;
  wire[0:0] quadInters_run_quadInters_run_or_46_nl;
  wire[0:0] quadInters_run_quadInters_run_or_48_nl;
  wire[31:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_mux_nl;
  wire[0:0] nor_74_nl;
  wire[0:0] quadInters_denom_dot_run_and_3_nl;
  wire[0:0] not_671_nl;
  wire[0:0] quad_hit_anything_mux_3_nl;
  wire[0:0] rec_quad_normal_z_not_nl;
  wire[0:0] rec_quad_normal_y_not_nl;
  wire[0:0] rec_quad_normal_x_not_nl;
  wire[27:0] quadInters_run_if_4_acc_nl;
  wire[28:0] nl_quadInters_run_if_4_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl;
  wire[57:0] quadInters_denom_dot_run_acc_2_nl;
  wire[58:0] nl_quadInters_denom_dot_run_acc_2_nl;
  wire[57:0] ac_math_ac_abs_58_58_xabs_xor_nl;
  wire[34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl;
  wire[35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_30_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_61_nl;
  wire[34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl;
  wire[35:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_62_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl;
  wire[0:0] quad_hit_anything_mux1h_58_nl;
  wire[0:0] setfacenorm_dot_run_and_1_nl;
  wire[22:0] quadInters_sub_run_acc_1_nl;
  wire[23:0] nl_quadInters_sub_run_acc_1_nl;
  wire[22:0] quadInters_sub_run_acc_2_nl;
  wire[23:0] nl_quadInters_sub_run_acc_2_nl;
  wire[22:0] quadInters_sub_run_acc_nl;
  wire[23:0] nl_quadInters_sub_run_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_73_nl;
  wire[34:0] quadInters_run_if_2_acc_nl;
  wire[35:0] nl_quadInters_run_if_2_acc_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl;
  wire[34:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_nl;
  wire[0:0] operator_35_true_mux_172_nl;
  wire[19:0] quadInters_run_mux_596_nl;
  wire[0:0] quadInters_run_and_2_nl;
  wire[19:0] quadInters_run_mux_595_nl;
  wire[0:0] quadInters_run_and_1_nl;
  wire[19:0] quadInters_run_mux_594_nl;
  wire[0:0] quadInters_run_and_nl;
  wire[47:0] quadInters_run_oif_acc_nl;
  wire[49:0] nl_quadInters_run_oif_acc_nl;
  wire[25:0] setfacenorm_negate_run_acc_2_nl;
  wire[26:0] nl_setfacenorm_negate_run_acc_2_nl;
  wire[25:0] setfacenorm_negate_run_acc_1_nl;
  wire[26:0] nl_setfacenorm_negate_run_acc_1_nl;
  wire[25:0] setfacenorm_negate_run_acc_nl;
  wire[26:0] nl_setfacenorm_negate_run_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_56_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_11_nl;
  wire[38:0] operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[39:0] nl_operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl;
  wire[38:0] operator_38_15_true_AC_TRN_AC_WRAP_acc_nl;
  wire[39:0] nl_operator_38_15_true_AC_TRN_AC_WRAP_acc_nl;
  wire[61:0] quadInters_beta_dot_run_acc_nl;
  wire[62:0] nl_quadInters_beta_dot_run_acc_nl;
  wire[61:0] quadInters_beta_dot_run_acc_2_nl;
  wire[62:0] nl_quadInters_beta_dot_run_acc_2_nl;
  wire[61:0] quadInters_alpha_dot_run_acc_nl;
  wire[62:0] nl_quadInters_alpha_dot_run_acc_nl;
  wire[61:0] quadInters_alpha_dot_run_acc_2_nl;
  wire[62:0] nl_quadInters_alpha_dot_run_acc_2_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_72_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_71_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_70_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_69_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_68_nl;
  wire[57:0] ac_math_ac_abs_58_58_xabs_acc_nl;
  wire[58:0] nl_ac_math_ac_abs_58_58_xabs_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_46_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_29_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_59_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_28_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_57_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_27_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_55_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_9_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_19_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_8_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_57_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_58_nl;
  wire[59:0] setfacenorm_dot_run_acc_nl;
  wire[60:0] nl_setfacenorm_dot_run_acc_nl;
  wire[21:0] quadInters_run_acc_6_nl;
  wire[22:0] nl_quadInters_run_acc_6_nl;
  wire[21:0] quadInters_run_acc_5_nl;
  wire[22:0] nl_quadInters_run_acc_5_nl;
  wire[20:0] ac_math_ac_abs_21_21_1_xabs_acc_nl;
  wire[21:0] nl_ac_math_ac_abs_21_21_1_xabs_acc_nl;
  wire[21:0] quadInters_run_acc_4_nl;
  wire[22:0] nl_quadInters_run_acc_4_nl;
  wire[20:0] ac_math_ac_abs_21_21_xabs_acc_nl;
  wire[21:0] nl_ac_math_ac_abs_21_21_xabs_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_77_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_76_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_75_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_74_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_54_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_53_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_52_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_55_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_34_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_33_nl;
  wire[59:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl;
  wire[60:0] nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_o000000;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_mux_nl;
  wire[47:0] quadInters_qnorm_rorig_run_acc_nl;
  wire[49:0] nl_quadInters_qnorm_rorig_run_acc_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_38_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_37_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_36_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_35_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_64_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_63_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_62_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_44_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_43_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_42_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_24_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_49_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_47_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_80_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_3_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_81_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_2_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_82_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_1_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_83_nl;
  wire[34:0] quadInters_run_if_1_acc_nl;
  wire[35:0] nl_quadInters_run_if_1_acc_nl;
  wire[60:0] acc_nl;
  wire[61:0] nl_acc_nl;
  wire[59:0] quadInters_cross_v_run_mux_2_nl;
  wire[56:0] quadInters_cross_v_run_mul_6_nl;
  wire[0:0] quadInters_cross_v_run_or_1_nl;
  wire[59:0] quadInters_cross_v_run_mux_3_nl;
  wire[56:0] quadInters_cross_v_run_mul_7_nl;
  wire[14:0] for_for_and_2_nl;
  wire[4:0] for_mux_25_nl;
  wire[0:0] for_or_11_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_21_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_131_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_132_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_82_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_83_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_84_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_133_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_85_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_123_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_124_nl;
  wire[34:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_125_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_86_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_126_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_87_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_127_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_128_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_129_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_88_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_89_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_130_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_131_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_132_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_133_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_90_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_91_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_134_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_135_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_136_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_137_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_92_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_93_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_138_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_139_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_94_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_95_nl;
  wire[32:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_140_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_14_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_134_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_15_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_96_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_97_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_16_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_22_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_141_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_142_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_23_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_135_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_98_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_99_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_136_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_24_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_143_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_144_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_100_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_101_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_145_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_146_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_147_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_102_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_103_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_2_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_49_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_50_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_148_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_104_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_149_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_25_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_150_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_151_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_152_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_105_nl;
  wire[33:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_153_nl;
  wire[0:0] div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_26_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [225:0] nl_IntersecLoop_hit_rec_quad_out_rsci_inst_rec_quad_out_rsci_idat;
  assign nl_IntersecLoop_hit_rec_quad_out_rsci_inst_rec_quad_out_rsci_idat = {rec_quad_out_rsci_idat_225_199
      , rec_quad_out_rsci_idat_198_172 , rec_quad_out_rsci_idat_171_145 , rec_quad_out_rsci_idat_144_142
      , rec_quad_out_rsci_idat_141 , rec_quad_out_rsci_idat_140_115 , rec_quad_out_rsci_idat_114_89
      , rec_quad_out_rsci_idat_88_63 , rec_quad_out_rsci_idat_62_43 , rec_quad_out_rsci_idat_42
      , rec_quad_out_rsci_idat_41_22 , rec_quad_out_rsci_idat_21 , rec_quad_out_rsci_idat_20_1
      , rec_quad_out_rsci_idat_0};
  wire [46:0] nl_IntersecLoop_hit_closest_so_far_out_rsci_inst_closest_so_far_out_rsci_idat;
  assign nl_IntersecLoop_hit_closest_so_far_out_rsci_inst_closest_so_far_out_rsci_idat
      = {closest_so_far_out_rsci_idat_46 , closest_so_far_out_rsci_idat_45 , closest_so_far_out_rsci_idat_44
      , closest_so_far_out_rsci_idat_43 , closest_so_far_out_rsci_idat_42 , closest_so_far_out_rsci_idat_41
      , closest_so_far_out_rsci_idat_40 , closest_so_far_out_rsci_idat_39 , closest_so_far_out_rsci_idat_38
      , closest_so_far_out_rsci_idat_37 , closest_so_far_out_rsci_idat_36 , closest_so_far_out_rsci_idat_35
      , closest_so_far_out_rsci_idat_34 , closest_so_far_out_rsci_idat_33 , closest_so_far_out_rsci_idat_32
      , closest_so_far_out_rsci_idat_31 , closest_so_far_out_rsci_idat_30 , closest_so_far_out_rsci_idat_29
      , closest_so_far_out_rsci_idat_28 , closest_so_far_out_rsci_idat_27 , closest_so_far_out_rsci_idat_26
      , closest_so_far_out_rsci_idat_25 , closest_so_far_out_rsci_idat_24 , closest_so_far_out_rsci_idat_23
      , closest_so_far_out_rsci_idat_22 , closest_so_far_out_rsci_idat_21 , closest_so_far_out_rsci_idat_20
      , closest_so_far_out_rsci_idat_19 , closest_so_far_out_rsci_idat_18 , closest_so_far_out_rsci_idat_17
      , closest_so_far_out_rsci_idat_16 , closest_so_far_out_rsci_idat_15 , closest_so_far_out_rsci_idat_14
      , closest_so_far_out_rsci_idat_13 , closest_so_far_out_rsci_idat_12 , closest_so_far_out_rsci_idat_11
      , closest_so_far_out_rsci_idat_10 , closest_so_far_out_rsci_idat_9 , closest_so_far_out_rsci_idat_8
      , closest_so_far_out_rsci_idat_7 , closest_so_far_out_rsci_idat_6 , closest_so_far_out_rsci_idat_5
      , closest_so_far_out_rsci_idat_4 , closest_so_far_out_rsci_idat_3 , closest_so_far_out_rsci_idat_2
      , closest_so_far_out_rsci_idat_1 , closest_so_far_out_rsci_idat_0};
  IntersecLoop_hit_quads_rsci IntersecLoop_hit_quads_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsc_dat(quads_rsc_dat),
      .quads_rsc_vld(quads_rsc_vld),
      .quads_rsc_rdy(quads_rsc_rdy),
      .hit_wen(hit_wen),
      .quads_rsci_oswt(reg_quads_rsci_irdy_hit_psct_cse),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .quads_rsci_idat_mxwt(quads_rsci_idat_mxwt)
    );
  IntersecLoop_hit_ray_temp_in_rsci IntersecLoop_hit_ray_temp_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_temp_in_rsc_dat(ray_temp_in_rsc_dat),
      .ray_temp_in_rsc_vld(ray_temp_in_rsc_vld),
      .ray_temp_in_rsc_rdy(ray_temp_in_rsc_rdy),
      .hit_wen(hit_wen),
      .ray_temp_in_rsci_oswt(reg_quad_max_in_rsci_irdy_hit_psct_cse),
      .ray_temp_in_rsci_wen_comp(ray_temp_in_rsci_wen_comp),
      .ray_temp_in_rsci_idat_mxwt(ray_temp_in_rsci_idat_mxwt)
    );
  IntersecLoop_hit_quad_max_in_rsci IntersecLoop_hit_quad_max_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quad_max_in_rsc_dat(quad_max_in_rsc_dat),
      .quad_max_in_rsc_vld(quad_max_in_rsc_vld),
      .quad_max_in_rsc_rdy(quad_max_in_rsc_rdy),
      .hit_wen(hit_wen),
      .quad_max_in_rsci_oswt(reg_quad_max_in_rsci_irdy_hit_psct_cse),
      .quad_max_in_rsci_wen_comp(quad_max_in_rsci_wen_comp),
      .quad_max_in_rsci_idat_mxwt(quad_max_in_rsci_idat_mxwt)
    );
  IntersecLoop_hit_quad_hit_anything_out_rsci IntersecLoop_hit_quad_hit_anything_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_out_rsc_dat(quad_hit_anything_out_rsc_dat),
      .quad_hit_anything_out_rsc_vld(quad_hit_anything_out_rsc_vld),
      .quad_hit_anything_out_rsc_rdy(quad_hit_anything_out_rsc_rdy),
      .hit_wen(hit_wen),
      .quad_hit_anything_out_rsci_oswt(reg_closest_so_far_out_rsci_ivld_hit_psct_cse),
      .quad_hit_anything_out_rsci_wen_comp(quad_hit_anything_out_rsci_wen_comp),
      .quad_hit_anything_out_rsci_idat(quad_hit_anything_out_rsci_idat)
    );
  IntersecLoop_hit_rec_quad_out_rsci IntersecLoop_hit_rec_quad_out_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_out_rsc_dat(rec_quad_out_rsc_dat),
      .rec_quad_out_rsc_vld(rec_quad_out_rsc_vld),
      .rec_quad_out_rsc_rdy(rec_quad_out_rsc_rdy),
      .hit_wen(hit_wen),
      .rec_quad_out_rsci_oswt(reg_closest_so_far_out_rsci_ivld_hit_psct_cse),
      .rec_quad_out_rsci_wen_comp(rec_quad_out_rsci_wen_comp),
      .rec_quad_out_rsci_idat(nl_IntersecLoop_hit_rec_quad_out_rsci_inst_rec_quad_out_rsci_idat[225:0])
    );
  IntersecLoop_hit_closest_so_far_out_rsci IntersecLoop_hit_closest_so_far_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_out_rsc_dat(closest_so_far_out_rsc_dat),
      .closest_so_far_out_rsc_vld(closest_so_far_out_rsc_vld),
      .closest_so_far_out_rsc_rdy(closest_so_far_out_rsc_rdy),
      .hit_wen(hit_wen),
      .closest_so_far_out_rsci_oswt(reg_closest_so_far_out_rsci_ivld_hit_psct_cse),
      .closest_so_far_out_rsci_wen_comp(closest_so_far_out_rsci_wen_comp),
      .closest_so_far_out_rsci_idat(nl_IntersecLoop_hit_closest_so_far_out_rsci_inst_closest_so_far_out_rsci_idat[46:0])
    );
  IntersecLoop_hit_wait_dp IntersecLoop_hit_wait_dp_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ensig_cgo_iro(ensig_cgo_mx0),
      .mult_run_mul_cmp_en(mult_run_mul_cmp_en),
      .mult_run_mul_cmp_z(mult_run_mul_cmp_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_z(quadInters_qnorm_rorig_run_mul_1_cmp_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_1_z(quadInters_qnorm_rorig_run_mul_1_cmp_1_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_2_z(quadInters_qnorm_rorig_run_mul_1_cmp_2_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_3_z(quadInters_qnorm_rorig_run_mul_1_cmp_3_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_4_z(quadInters_qnorm_rorig_run_mul_1_cmp_4_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_5_z(quadInters_qnorm_rorig_run_mul_1_cmp_5_z),
      .quadInters_denom_dot_run_mul_2_cmp_z(quadInters_denom_dot_run_mul_2_cmp_z),
      .quadInters_denom_dot_run_mul_2_cmp_1_z(quadInters_denom_dot_run_mul_2_cmp_1_z),
      .quadInters_denom_dot_run_mul_1_cmp_z(quadInters_denom_dot_run_mul_1_cmp_z),
      .hit_wen(hit_wen),
      .ensig_cgo(ensig_cgo),
      .mult_run_mul_cmp_z_oreg(mult_run_mul_cmp_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg),
      .quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg(quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg),
      .quadInters_denom_dot_run_mul_2_cmp_z_oreg(quadInters_denom_dot_run_mul_2_cmp_z_oreg),
      .quadInters_denom_dot_run_mul_2_cmp_1_z_oreg(quadInters_denom_dot_run_mul_2_cmp_1_z_oreg),
      .quadInters_denom_dot_run_mul_1_cmp_z_oreg(quadInters_denom_dot_run_mul_1_cmp_z_oreg)
    );
  IntersecLoop_hit_staller IntersecLoop_hit_staller_inst (
      .hit_wen(hit_wen),
      .quads_rsci_wen_comp(quads_rsci_wen_comp),
      .ray_temp_in_rsci_wen_comp(ray_temp_in_rsci_wen_comp),
      .quad_max_in_rsci_wen_comp(quad_max_in_rsci_wen_comp),
      .quad_hit_anything_out_rsci_wen_comp(quad_hit_anything_out_rsci_wen_comp),
      .rec_quad_out_rsci_wen_comp(rec_quad_out_rsci_wen_comp),
      .closest_so_far_out_rsci_wen_comp(closest_so_far_out_rsci_wen_comp)
    );
  IntersecLoop_hit_hit_fsm IntersecLoop_hit_hit_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .hit_wen(hit_wen),
      .fsm_output(fsm_output),
      .for_C_3_tr0(for_nor_tmp)
    );
  assign closest_so_far_out_and_cse = hit_wen & (fsm_output[5]) & for_nor_tmp;
  assign closest_so_far_and_cse = hit_wen & (or_tmp_328 | (fsm_output[5]));
  assign closest_so_far_and_47_cse = closest_so_far_and_cse & (for_stage_0_8 | (~
      (fsm_output[5])));
  assign rec_quad_color_b_and_cse = hit_wen & (((~ quadInters_run_if_5_quadInters_run_if_5_or_2_tmp)
      & (~(quadInters_run_lor_lpi_2_dfm_1 | quadInters_run_land_lpi_2_dfm_8)) & (~
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7) & for_stage_0_9 &
      (fsm_output[2])) | or_tmp_328);
  assign rec_quad_normal_z_and_cse = hit_wen & (or_tmp_480 | or_tmp_481);
  assign rec_quad_hit_loc_z_and_cse = hit_wen & ((for_hitWorld_lpi_2_dfm_2 & for_stage_0_9
      & (fsm_output[3])) | or_tmp_490);
  assign add_run_and_3_cse = hit_wen & (~(quadInters_run_land_lpi_2_dfm_st_7 | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6
      | (~ for_stage_0_8))) & (fsm_output[3]);
  assign rec_quad_mat_and_1_rgt = for_stage_0_8 & (fsm_output[5]);
  assign ac_math_ac_abs_21_21_1_xabs_and_1_cse = for_stage_0_9 & (fsm_output[2]);
  assign or_cse = (fsm_output[3:2]!=2'b00);
  assign and_2744_cse = ((or_cse & for_stage_0_9) | (fsm_output[0])) & hit_wen;
  assign quadInters_run_oelse_and_1_cse = hit_wen & (fsm_output[5]);
  assign and_2754_cse = (~((~(for_stage_0_9 & for_hitWorld_lpi_2_dfm_2 & (~ operator_33_true_asn_1_itm_8)))
      & (fsm_output[3]))) & (~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[2])))
      & hit_wen;
  assign and_2778_cse = (~((~(for_stage_0_9 & (~ quadInters_run_lor_lpi_2_dfm_1)
      & (~ (quadInters_alpha_dot_run_acc_itm_61_24[37])) & (~(operator_33_true_asn_1_itm_8
      | quadInters_run_land_lpi_2_dfm_8)) & (~(quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7
      | operator_38_15_true_AC_TRN_AC_WRAP_acc_itm_38)) & (~((quadInters_beta_dot_run_acc_itm_61_24[37])
      | operator_38_15_true_AC_TRN_AC_WRAP_1_acc_itm_38)))) & (fsm_output[2]))) &
      (fsm_output[5:3]==3'b000) & hit_wen;
  assign quadInters_run_t_trunc_mux_47_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_46,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46,
      fsm_output[5]);
  assign quadInters_run_t_trunc_mux_48_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_45,
      quadInters_run_t_trunc_lpi_2_dfm_45_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_49_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_44,
      quadInters_run_t_trunc_lpi_2_dfm_44_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_50_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_43,
      quadInters_run_t_trunc_lpi_2_dfm_43_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_51_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_42,
      quadInters_run_t_trunc_lpi_2_dfm_42_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_52_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_41,
      quadInters_run_t_trunc_lpi_2_dfm_41_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_53_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_40,
      quadInters_run_t_trunc_lpi_2_dfm_40_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_54_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_39,
      quadInters_run_t_trunc_lpi_2_dfm_39_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_55_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_38,
      quadInters_run_t_trunc_lpi_2_dfm_38_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_56_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_37,
      quadInters_run_t_trunc_lpi_2_dfm_37_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_57_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_36,
      quadInters_run_t_trunc_lpi_2_dfm_36_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_58_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_35,
      quadInters_run_t_trunc_lpi_2_dfm_35_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_59_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_34,
      quadInters_run_t_trunc_lpi_2_dfm_34_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_60_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_33,
      quadInters_run_t_trunc_lpi_2_dfm_33_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_61_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_32,
      quadInters_run_t_trunc_lpi_2_dfm_32_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_62_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_31,
      quadInters_run_t_trunc_lpi_2_dfm_31_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_63_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_30,
      quadInters_run_t_trunc_lpi_2_dfm_30_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_64_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_29,
      quadInters_run_t_trunc_lpi_2_dfm_29_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_65_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_28,
      quadInters_run_t_trunc_lpi_2_dfm_28_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_66_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_27,
      quadInters_run_t_trunc_lpi_2_dfm_27_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_67_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_26,
      quadInters_run_t_trunc_lpi_2_dfm_26_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_68_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_25,
      quadInters_run_t_trunc_lpi_2_dfm_25_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_69_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_24,
      quadInters_run_t_trunc_lpi_2_dfm_24_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_70_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_23,
      quadInters_run_t_trunc_lpi_2_dfm_23_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_71_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_22,
      quadInters_run_t_trunc_lpi_2_dfm_22_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_72_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_21,
      quadInters_run_t_trunc_lpi_2_dfm_21_1, fsm_output[5]);
  assign quadInters_run_t_trunc_mux_73_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_20,
      quadInters_run_t_trunc_lpi_2_dfm_20_1, fsm_output[5]);
  assign quadInters_run_quadInters_run_or_10_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_74_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_19,
      (quadInters_run_quadInters_run_or_10_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_12_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_75_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_18,
      (quadInters_run_quadInters_run_or_12_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_14_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_76_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_17,
      (quadInters_run_quadInters_run_or_14_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_16_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_77_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_16,
      (quadInters_run_quadInters_run_or_16_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_18_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_78_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_15,
      (quadInters_run_quadInters_run_or_18_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_20_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_79_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_14,
      (quadInters_run_quadInters_run_or_20_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_22_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_80_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_13,
      (quadInters_run_quadInters_run_or_22_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_24_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_81_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_12,
      (quadInters_run_quadInters_run_or_24_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_26_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_82_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_11,
      (quadInters_run_quadInters_run_or_26_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_28_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_83_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_10,
      (quadInters_run_quadInters_run_or_28_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_30_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_9
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_84_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_9,
      (quadInters_run_quadInters_run_or_30_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_32_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_8
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_85_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_8,
      (quadInters_run_quadInters_run_or_32_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_34_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_7
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_86_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_7,
      (quadInters_run_quadInters_run_or_34_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_36_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_6
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_87_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_6,
      (quadInters_run_quadInters_run_or_36_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_38_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_5
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_88_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_5,
      (quadInters_run_quadInters_run_or_38_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_40_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_4
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_89_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_4,
      (quadInters_run_quadInters_run_or_40_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_42_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_90_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_3,
      (quadInters_run_quadInters_run_or_42_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_44_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_91_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_2,
      (quadInters_run_quadInters_run_or_44_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_46_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_92_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_1,
      (quadInters_run_quadInters_run_or_46_nl), fsm_output[5]);
  assign quadInters_run_quadInters_run_or_48_nl = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_mux_93_cse = MUX_s_1_2_2(quadInters_run_t_trunc_lpi_2_dfm_1_0,
      (quadInters_run_quadInters_run_or_48_nl), fsm_output[5]);
  assign quadInters_denom_dot_run_and_4_rgt = (~ quadInters_run_land_lpi_2_dfm) &
      (fsm_output[5]);
  assign quadInters_denom_dot_run_and_5_rgt = quadInters_run_land_lpi_2_dfm & (fsm_output[5]);
  assign nor_74_nl = ~(quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs | (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_mux_nl
      = MUX_v_32_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0[31:0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[31:0]),
      nor_74_nl);
  assign quadInters_denom_dot_run_and_3_nl = (~(quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs
      | (~ quadInters_run_if_1_acc_itm_34))) & (fsm_output[3]);
  assign quadInters_denom_dot_run_mux1h_5_rgt = MUX1HOT_v_34_4_2(({{32{quadInters_run_if_1_exs_mx1w0_1_0[1]}},
      quadInters_run_if_1_exs_mx1w0_1_0}), ({2'b00 , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qelse_mux_nl)}),
      (quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0[57:24]), quadInters_denom_dot_run_ac_fixed_cctor_sva_57_24,
      {(quadInters_denom_dot_run_and_3_nl) , (fsm_output[4]) , quadInters_denom_dot_run_and_4_rgt
      , quadInters_denom_dot_run_and_5_rgt});
  assign or_343_cse = (((for_i_5_0_sva_4_0) == (operator_11_false_acc_sdt_sva_1[4:0]))
      & (operator_11_false_acc_sdt_sva_1[11:5]==7'b0000000)) | (z_out_1[5]);
  assign and_1706_cse = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
      & (~ operator_33_true_asn_1_itm_9) & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st
      & (fsm_output[3]);
  assign and_2828_cse = (and_1706_cse | (fsm_output[6]) | (fsm_output[0]) | (fsm_output[1]))
      & hit_wen;
  assign and_2843_cse = (~(operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm
      | quadInters_run_land_lpi_2_dfm_9)) & (~(quadInters_run_lor_3_lpi_2_dfm_1 |
      quadInters_run_lor_lpi_2_dfm_2)) & (fsm_output[3]) & (~ operator_33_true_asn_1_itm_9)
      & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
      & hit_wen;
  assign quadInters_run_oelse_and_2_cse = hit_wen & (~((fsm_output[4]) | (fsm_output[2])));
  assign operator_35_true_and_57_cse = (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4)
      & (fsm_output[4]);
  assign operator_35_true_and_58_cse = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4
      & (fsm_output[4]);
  assign operator_35_true_and_30_rgt = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3
      & (fsm_output[5]);
  assign operator_35_true_and_31_rgt = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3)
      & (fsm_output[5]);
  assign operator_35_true_and_32_rgt = (~(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3))
      & (fsm_output[5]);
  assign operator_35_true_and_59_cse = hit_wen & (~ or_cse);
  assign for_and_1_cse = hit_wen & ((fsm_output[5]) | (fsm_output[1]));
  assign operator_35_true_and_100_cse = hit_wen & (~((~ for_stage_0_5) | quadInters_run_land_lpi_2_dfm_st_4
      | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3 | (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3)))
      & (fsm_output[5]);
  assign operator_35_true_and_282_cse = and_dcpl_238 & (fsm_output[5]);
  assign operator_35_true_and_135_cse = hit_wen & (((quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2
      | quadInters_run_land_lpi_2_dfm_st_3 | (~(for_stage_0_4 & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2)))
      & for_stage_0_5 & (~ quadInters_run_land_lpi_2_dfm_st_4) & (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3)
      & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3)
      | and_dcpl_238) & (fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_cse
      = hit_wen & (~ or_dcpl_79);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_3_cse
      = hit_wen & (~ (fsm_output[4]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_6_rgt
      = (~(quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs | (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0[34])))
      & (fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_m1c
      = (fsm_output[5:3]!=3'b000);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_11_rgt
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1,
      z_out_2, fsm_output[5]);
  assign or_1462_cse = (fsm_output[5:4]!=2'b00);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_1_cse
      = quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs & (fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_or_rgt
      = or_cse | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_1_cse;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_rgt
      = (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs) & (fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_5_cse
      = hit_wen & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_or_rgt);
  assign operator_35_true_and_16_rgt = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3
      & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3
      & (fsm_output[5]);
  assign operator_35_true_and_185_cse = hit_wen & (~(or_cse | ((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3)
      & (fsm_output[5]))));
  assign nl_quadInters_sub_run_acc_1_nl = (add_run_ac_fixed_cctor_1_74_43_sva_mx1w0[31:9])
      - conv_s2u_12_23(quads_crt_sva_7_110_0[23:12]);
  assign quadInters_sub_run_acc_1_nl = nl_quadInters_sub_run_acc_1_nl[22:0];
  assign quadInters_sub_run_mux_rgt = MUX_v_23_2_2(({2'b00 , (add_run_ac_fixed_cctor_1_74_43_sva[20:0])}),
      (quadInters_sub_run_acc_1_nl), fsm_output[3]);
  assign and_2862_cse = ((fsm_output[5]) | (fsm_output[3])) & hit_wen;
  assign nl_quadInters_sub_run_acc_2_nl = (add_run_ac_fixed_cctor_2_74_43_sva_mx1w0[31:9])
      - conv_s2u_12_23(quads_crt_sva_7_110_0[35:24]);
  assign quadInters_sub_run_acc_2_nl = nl_quadInters_sub_run_acc_2_nl[22:0];
  assign quadInters_sub_run_mux_1_rgt = MUX_v_23_2_2(({2'b00 , (add_run_ac_fixed_cctor_2_74_43_sva[20:0])}),
      (quadInters_sub_run_acc_2_nl), fsm_output[3]);
  assign nl_quadInters_sub_run_acc_nl = (add_run_ac_fixed_cctor_74_43_sva_mx1w0[31:9])
      - conv_s2u_12_23(quads_crt_sva_7_110_0[11:0]);
  assign quadInters_sub_run_acc_nl = nl_quadInters_sub_run_acc_nl[22:0];
  assign quadInters_sub_run_mux_2_rgt = MUX_v_23_2_2(({2'b00 , (add_run_ac_fixed_cctor_74_43_sva[20:0])}),
      (quadInters_sub_run_acc_nl), fsm_output[3]);
  assign and_2865_cse = (~ (fsm_output[3])) & hit_wen;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_73_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_73_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_73_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_74_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_and_rgt
      = ~(quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs | quadInters_run_mux_593_tmp_33
      | (fsm_output[4]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_cse
      = hit_wen & and_454_cse;
  assign and_454_cse = (~(quadInters_run_land_lpi_2_dfm_st_5 | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_4))
      & for_stage_0_6;
  assign ensig_cgo_mx0 = (and_dcpl_195 & or_dcpl_79) | ((and_dcpl_195 | and_454_cse)
      & (fsm_output[5])) | ((and_dcpl_54 | and_dcpl_195) & (fsm_output[2]));
  assign quad_hit_anything_sva_dfm_mx0w0 = quad_hit_anything_sva | for_hitWorld_lpi_2_dfm_3;
  assign quadInters_run_quadInters_run_quadInters_run_nor_6_mx0w1 = ~((~((reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg[0])
      | quadInters_run_acc_6_itm_21)) | quadInters_run_lor_3_lpi_2_dfm | quadInters_run_lor_lpi_2_dfm_1
      | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 | quadInters_run_land_lpi_2_dfm_8);
  assign quadInters_run_and_2_nl = quadInters_run_acc_6_itm_21 & (~ quadInters_run_lor_3_lpi_2_dfm);
  assign quadInters_run_mux_596_nl = MUX_v_20_2_2((reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg[20:1]),
      ({{19{div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}},
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}),
      quadInters_run_and_2_nl);
  assign quadInters_run_quadInters_run_and_6_mx0w2 = (quadInters_run_mux_596_nl)
      & (signext_20_1(~ quadInters_run_lor_3_lpi_2_dfm)) & (signext_20_1(~ quadInters_run_lor_lpi_2_dfm_1))
      & (signext_20_1(~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7))
      & (signext_20_1(~ quadInters_run_land_lpi_2_dfm_8));
  assign quadInters_run_quadInters_run_quadInters_run_nor_5_mx0w1 = ~((~((reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg[0])
      | quadInters_run_acc_5_itm_21)) | quadInters_run_lor_3_lpi_2_dfm | quadInters_run_lor_lpi_2_dfm_1
      | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 | quadInters_run_land_lpi_2_dfm_8);
  assign quadInters_run_and_1_nl = quadInters_run_acc_5_itm_21 & (~ quadInters_run_lor_3_lpi_2_dfm);
  assign quadInters_run_mux_595_nl = MUX_v_20_2_2((reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg[20:1]),
      ({{19{div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}},
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}),
      quadInters_run_and_1_nl);
  assign quadInters_run_quadInters_run_and_4_mx0w2 = (quadInters_run_mux_595_nl)
      & (signext_20_1(~ quadInters_run_lor_3_lpi_2_dfm)) & (signext_20_1(~ quadInters_run_lor_lpi_2_dfm_1))
      & (signext_20_1(~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7))
      & (signext_20_1(~ quadInters_run_land_lpi_2_dfm_8));
  assign quadInters_run_quadInters_run_quadInters_run_nor_mx0w1 = ~((~((reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg[0])
      | quadInters_run_acc_4_itm_21)) | quadInters_run_lor_3_lpi_2_dfm | quadInters_run_lor_lpi_2_dfm_1
      | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 | quadInters_run_land_lpi_2_dfm_8);
  assign quadInters_run_and_nl = quadInters_run_acc_4_itm_21 & (~ quadInters_run_lor_3_lpi_2_dfm);
  assign quadInters_run_mux_594_nl = MUX_v_20_2_2((reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg[20:1]),
      ({{19{div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}},
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm}),
      quadInters_run_and_nl);
  assign quadInters_run_quadInters_run_and_2_mx0w2 = (quadInters_run_mux_594_nl)
      & (signext_20_1(~ quadInters_run_lor_3_lpi_2_dfm)) & (signext_20_1(~ quadInters_run_lor_lpi_2_dfm_1))
      & (signext_20_1(~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7))
      & (signext_20_1(~ quadInters_run_land_lpi_2_dfm_8));
  assign nl_add_run_ac_fixed_cctor_2_74_43_sva_mx1w0 = conv_s2u_21_32(ray_temp_in_crt_sva[62:42])
      + (mult_run_asn_2_itm_1_74_30[44:13]);
  assign add_run_ac_fixed_cctor_2_74_43_sva_mx1w0 = nl_add_run_ac_fixed_cctor_2_74_43_sva_mx1w0[31:0];
  assign nl_add_run_ac_fixed_cctor_1_74_43_sva_mx1w0 = conv_s2u_21_32(ray_temp_in_crt_sva[41:21])
      + mult_run_asn_1_itm_74_43;
  assign add_run_ac_fixed_cctor_1_74_43_sva_mx1w0 = nl_add_run_ac_fixed_cctor_1_74_43_sva_mx1w0[31:0];
  assign nl_add_run_ac_fixed_cctor_74_43_sva_mx1w0 = conv_s2u_21_32(ray_temp_in_crt_sva[20:0])
      + (mult_run_mul_cmp_z_oreg[44:13]);
  assign add_run_ac_fixed_cctor_74_43_sva_mx1w0 = nl_add_run_ac_fixed_cctor_74_43_sva_mx1w0[31:0];
  assign nl_quadInters_run_oif_acc_nl = conv_s2u_47_48({closest_so_far_sva_46 , closest_so_far_sva_45
      , closest_so_far_sva_44 , closest_so_far_sva_43 , closest_so_far_sva_42 , closest_so_far_sva_41
      , closest_so_far_sva_40 , closest_so_far_sva_39 , closest_so_far_sva_38 , closest_so_far_sva_37
      , closest_so_far_sva_36 , closest_so_far_sva_35 , closest_so_far_sva_34 , closest_so_far_sva_33
      , closest_so_far_sva_32 , closest_so_far_sva_31 , closest_so_far_sva_30 , closest_so_far_sva_29
      , closest_so_far_sva_28 , closest_so_far_sva_27 , closest_so_far_sva_26 , closest_so_far_sva_25
      , closest_so_far_sva_24 , closest_so_far_sva_23 , closest_so_far_sva_22 , closest_so_far_sva_21
      , closest_so_far_sva_20 , closest_so_far_sva_19 , closest_so_far_sva_18 , closest_so_far_sva_17
      , closest_so_far_sva_16 , closest_so_far_sva_15 , closest_so_far_sva_14 , closest_so_far_sva_13
      , closest_so_far_sva_12 , closest_so_far_sva_11 , closest_so_far_sva_10 , closest_so_far_sva_9
      , closest_so_far_sva_8 , closest_so_far_sva_7 , closest_so_far_sva_6 , closest_so_far_sva_5
      , closest_so_far_sva_4 , closest_so_far_sva_3 , closest_so_far_sva_2 , closest_so_far_sva_1
      , closest_so_far_sva_0}) + conv_s2u_47_48({(~ quadInters_run_t_trunc_lpi_2_dfm_2_46)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_45) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_44)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_43) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_42)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_41) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_40)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_39) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_38)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_37) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_36)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_35) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_34)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_33) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_32)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_31) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_30)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_29) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_28)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_27) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_26)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_25) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_24)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_23) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_22)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_21) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_20)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_19) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_18)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_17) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_16)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_15) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_14)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_13) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_12)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_11) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_10)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_9) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_8)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_7) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_6)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_5) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_4)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_3) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_2)
      , (~ quadInters_run_t_trunc_lpi_2_dfm_2_1) , (~ quadInters_run_t_trunc_lpi_2_dfm_2_0)})
      + 48'b000000000000000000000000000000000000000000000001;
  assign quadInters_run_oif_acc_nl = nl_quadInters_run_oif_acc_nl[47:0];
  assign quadInters_run_lor_lpi_2_dfm_mx0w1 = (readslicef_48_1_47((quadInters_run_oif_acc_nl)))
      | operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_33_itm;
  assign quadInters_run_t_trunc_lpi_2_dfm_45_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_45
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_44_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_44
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_43_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_43
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_42_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_42
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_41_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_41
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_40_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_40
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_39_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_39
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_38_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_38
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_37_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_37
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_36_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_36
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_35_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_35
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_34_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_34
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_33_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_33
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_32_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_32
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_31_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_31
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_30_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_30
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_29_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_29
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_28_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_28
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_27_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_27
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_26_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_26
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_25_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_25
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_24_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_24
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_23_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_23
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_22_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_22
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_21_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_21
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_t_trunc_lpi_2_dfm_20_1 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_itm
      | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46;
  assign quadInters_run_if_1_exs_mx1w0_1_0 = MUX_v_2_2_2(2'b01, 2'b10, quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56[1]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0
      = conv_u2u_33_34(~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[32:0]))
      + 34'b0000000000000000000000000000000001;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0[33:0];
  assign nl_setfacenorm_negate_run_acc_2_nl =  -(quads_crt_sva_9_189_112[77:52]);
  assign setfacenorm_negate_run_acc_2_nl = nl_setfacenorm_negate_run_acc_2_nl[25:0];
  assign quadInters_setfacenorm_run_qr_z_lpi_2_dfm_4_mx1w0 = MUX1HOT_v_26_3_2((setfacenorm_negate_run_acc_2_nl),
      (quads_crt_sva_9_189_112[77:52]), quadInters_setfacenorm_run_qr_z_lpi_2, {quadInters_run_asn_69
      , quadInters_run_quadInters_run_nor_4_cse_1 , quadInters_run_asn_71});
  assign nl_setfacenorm_negate_run_acc_1_nl =  -(quads_crt_sva_9_189_112[51:26]);
  assign setfacenorm_negate_run_acc_1_nl = nl_setfacenorm_negate_run_acc_1_nl[25:0];
  assign quadInters_setfacenorm_run_qr_y_lpi_2_dfm_4_mx1w0 = MUX1HOT_v_26_3_2((setfacenorm_negate_run_acc_1_nl),
      (quads_crt_sva_9_189_112[51:26]), quadInters_setfacenorm_run_qr_y_lpi_2, {quadInters_run_asn_69
      , quadInters_run_quadInters_run_nor_4_cse_1 , quadInters_run_asn_71});
  assign nl_setfacenorm_negate_run_acc_nl =  -(quads_crt_sva_9_189_112[25:0]);
  assign setfacenorm_negate_run_acc_nl = nl_setfacenorm_negate_run_acc_nl[25:0];
  assign quadInters_setfacenorm_run_qr_x_lpi_2_dfm_4_mx1w0 = MUX1HOT_v_26_3_2((setfacenorm_negate_run_acc_nl),
      (quads_crt_sva_9_189_112[25:0]), quadInters_setfacenorm_run_qr_x_lpi_2, {quadInters_run_asn_69
      , quadInters_run_quadInters_run_nor_4_cse_1 , quadInters_run_asn_71});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx1
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      z_out_5[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx2
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx3
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      z_out_5[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_56_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1
      = ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_32_0
      , (ac_math_ac_abs_58_58_xabs_57_24_sva[0])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_56_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_57_lpi_2_dfm[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1[33:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0
      = (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm)
      + 34'b0000000000000000000000000000000001;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_11_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1[33:0])
      , (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[27])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_11_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_mx1w0
      = ~((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[33])
      ^ (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56[1]));
  assign nl_operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl = conv_s2s_38_39(~ quadInters_beta_dot_run_acc_itm_61_24)
      + 39'b000000000000000100000000000000000000001;
  assign operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl = nl_operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl[38:0];
  assign operator_38_15_true_AC_TRN_AC_WRAP_1_acc_itm_38 = readslicef_39_1_38((operator_38_15_true_AC_TRN_AC_WRAP_1_acc_nl));
  assign nl_operator_38_15_true_AC_TRN_AC_WRAP_acc_nl = conv_s2s_38_39(~ quadInters_alpha_dot_run_acc_itm_61_24)
      + 39'b000000000000000100000000000000000000001;
  assign operator_38_15_true_AC_TRN_AC_WRAP_acc_nl = nl_operator_38_15_true_AC_TRN_AC_WRAP_acc_nl[38:0];
  assign operator_38_15_true_AC_TRN_AC_WRAP_acc_itm_38 = readslicef_39_1_38((operator_38_15_true_AC_TRN_AC_WRAP_acc_nl));
  assign quadInters_run_if_5_quadInters_run_if_5_or_2_tmp = operator_38_15_true_AC_TRN_AC_WRAP_1_acc_itm_38
      | (quadInters_beta_dot_run_acc_itm_61_24[37]) | operator_38_15_true_AC_TRN_AC_WRAP_acc_itm_38
      | (quadInters_alpha_dot_run_acc_itm_61_24[37]);
  assign for_hitWorld_lpi_2_dfm_3 = ~(quadInters_run_if_5_quadInters_run_if_5_or_2_tmp
      | quadInters_run_lor_lpi_2_dfm_1 | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7
      | quadInters_run_land_lpi_2_dfm_8);
  assign nl_quadInters_beta_dot_run_acc_2_nl = quadInters_qnorm_rorig_run_mul_1_cmp_1_z_oreg
      + quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg;
  assign quadInters_beta_dot_run_acc_2_nl = nl_quadInters_beta_dot_run_acc_2_nl[61:0];
  assign nl_quadInters_beta_dot_run_acc_nl = (quadInters_beta_dot_run_acc_2_nl) +
      quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg;
  assign quadInters_beta_dot_run_acc_nl = nl_quadInters_beta_dot_run_acc_nl[61:0];
  assign quadInters_beta_dot_run_acc_itm_61_24 = readslicef_62_38_24((quadInters_beta_dot_run_acc_nl));
  assign nl_quadInters_alpha_dot_run_acc_2_nl = quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg
      + quadInters_qnorm_rorig_run_mul_1_cmp_3_z_oreg;
  assign quadInters_alpha_dot_run_acc_2_nl = nl_quadInters_alpha_dot_run_acc_2_nl[61:0];
  assign nl_quadInters_alpha_dot_run_acc_nl = (quadInters_alpha_dot_run_acc_2_nl)
      + quadInters_qnorm_rorig_run_mul_1_cmp_2_z_oreg;
  assign quadInters_alpha_dot_run_acc_nl = nl_quadInters_alpha_dot_run_acc_nl[61:0];
  assign quadInters_alpha_dot_run_acc_itm_61_24 = readslicef_62_38_24((quadInters_alpha_dot_run_acc_nl));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_72_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_72_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_72_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_73_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_74_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_71_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_71_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_71_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_72_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_70_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_70_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_70_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_71_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_69_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_69_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_69_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_70_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_68_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1
      = ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_32_0
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_68_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_69_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_73_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_72_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_71_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_70_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_69_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33);
  assign nl_ac_math_ac_abs_58_58_xabs_acc_nl = ac_math_ac_abs_58_58_xabs_xor_itm
      + conv_u2u_1_58(quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56[1]);
  assign ac_math_ac_abs_58_58_xabs_acc_nl = nl_ac_math_ac_abs_58_58_xabs_acc_nl[57:0];
  assign ac_math_ac_abs_58_58_xabs_acc_itm_57_24 = readslicef_58_34_24((ac_math_ac_abs_58_58_xabs_acc_nl));
  assign ac_math_ac_abs_58_58_xabs_57_24_sva_mx1 = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[33]);
  assign nl_operator_11_false_acc_sdt_sva_1 = conv_u2s_11_12(quad_max_sva) + 12'b111111111111;
  assign operator_11_false_acc_sdt_sva_1 = nl_operator_11_false_acc_sdt_sva_1[11:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_48_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_49_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[32:0])
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_48_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_46_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1
      = ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_32_0
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_46_nl)
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_50_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_49_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_48_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[33]);
  assign nl_quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0 = ac_math_ac_abs_58_58_xabs_xor_itm
      + ({quadInters_denom_dot_run_ac_fixed_cctor_sva_57_24 , quadInters_denom_dot_run_ac_fixed_cctor_sva_23_0});
  assign quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0 = nl_quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0[57:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_29_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_59_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1[33:0])
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_3_itm_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_29_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_59_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_28_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_57_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1[33:0])
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_4_itm_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_28_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_57_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_27_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (z_out_10[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_55_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      z_out_10[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1
      = ({(z_out_10[33:0]) , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_5_itm_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_27_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_55_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_9_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_19_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1[33:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22[1])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_9_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_19_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_8_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_11[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      z_out_11[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1
      = ({(z_out_11[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22[2])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_8_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_11_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx0_33_32
      = MUX_v_2_2_2(({1'b0 , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[32])}),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx2w0[33:32]),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_mx2
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_57_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_57_lpi_2_dfm[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_57_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_58_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_58_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_58_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_58_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_59_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[33:0];
  assign nl_setfacenorm_dot_run_acc_nl = setfacenorm_dot_run_acc_2_itm + quadInters_denom_dot_run_mul_1_cmp_z_oreg;
  assign setfacenorm_dot_run_acc_nl = nl_setfacenorm_dot_run_acc_nl[59:0];
  assign setfacenorm_dot_run_acc_itm_59 = readslicef_60_1_59((setfacenorm_dot_run_acc_nl));
  assign quadInters_run_quadInters_run_nor_4_cse_1 = ~((~ setfacenorm_dot_run_acc_itm_59)
      | quadInters_run_lor_3_lpi_2_dfm_1 | quadInters_run_lor_lpi_2_dfm_2 | quadInters_run_or_1_tmp_1);
  assign quadInters_run_or_1_tmp_1 = operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm
      | quadInters_run_land_lpi_2_dfm_9;
  assign nl_quadInters_run_acc_6_nl = conv_s2u_21_22(z_out_1) + 22'b1111111111111111111111;
  assign quadInters_run_acc_6_nl = nl_quadInters_run_acc_6_nl[21:0];
  assign quadInters_run_acc_6_itm_21 = readslicef_22_1_21((quadInters_run_acc_6_nl));
  assign nl_ac_math_ac_abs_21_21_1_xabs_acc_nl = conv_u2s_20_21(reg_ac_math_ac_abs_21_21_1_xabs_xor_ftd_1)
      + conv_u2s_1_21(reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg[20]);
  assign ac_math_ac_abs_21_21_1_xabs_acc_nl = nl_ac_math_ac_abs_21_21_1_xabs_acc_nl[20:0];
  assign nl_quadInters_run_acc_5_nl = conv_s2u_21_22(ac_math_ac_abs_21_21_1_xabs_acc_nl)
      + 22'b1111111111111111111111;
  assign quadInters_run_acc_5_nl = nl_quadInters_run_acc_5_nl[21:0];
  assign quadInters_run_acc_5_itm_21 = readslicef_22_1_21((quadInters_run_acc_5_nl));
  assign nl_ac_math_ac_abs_21_21_xabs_acc_nl = conv_u2s_20_21(reg_ac_math_ac_abs_21_21_xabs_xor_ftd_1)
      + conv_u2s_1_21(reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg[20]);
  assign ac_math_ac_abs_21_21_xabs_acc_nl = nl_ac_math_ac_abs_21_21_xabs_acc_nl[20:0];
  assign nl_quadInters_run_acc_4_nl = conv_s2u_21_22(ac_math_ac_abs_21_21_xabs_acc_nl)
      + 22'b1111111111111111111111;
  assign quadInters_run_acc_4_nl = nl_quadInters_run_acc_4_nl[21:0];
  assign quadInters_run_acc_4_itm_21 = readslicef_22_1_21((quadInters_run_acc_4_nl));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_77_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_77_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_77_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_76_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_76_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_76_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_77_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_75_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_75_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_75_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_76_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_74_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1
      = ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_32_0
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_74_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_75_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_77_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_76_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_75_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33);
  assign quadInters_run_rounded_denom_lpi_2_dfm_mx0_32_0 = MUX_v_33_2_2(({(quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56[0])
      , quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24}), ({{31{quadInters_run_if_1_exs_mx1w0_1_0[1]}},
      quadInters_run_if_1_exs_mx1w0_1_0}), quadInters_run_if_1_acc_itm_34);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_54_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_54_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_54_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_55_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_53_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_53_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_53_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_54_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_52_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (z_out_7[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0
      = ({(z_out_7[32:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_52_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_52_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_53_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_55_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_55_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_55_nl)
      , (ac_math_ac_abs_58_58_xabs_57_24_sva_mx1[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_55_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_54_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_53_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      z_out_7[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_52_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_34_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_34_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_34_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_35_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_33_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (z_out_11[34]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1
      = (z_out_11[33:0]) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_33_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_34_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_35_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_34_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      z_out_11[34]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_13_cse
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_9[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_12_cse
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_10[34]));
  assign quadInters_run_asn_69 = ~(setfacenorm_dot_run_acc_itm_59 | quadInters_run_lor_3_lpi_2_dfm_1
      | quadInters_run_lor_lpi_2_dfm_2 | quadInters_run_or_1_tmp_1);
  assign quadInters_run_asn_71 = quadInters_run_lor_3_lpi_2_dfm_1 | quadInters_run_lor_lpi_2_dfm_2
      | quadInters_run_or_1_tmp_1;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_qelse_conc_itm_33
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (z_out_6[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1
      = ({(z_out_6[32:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_60_lpi_2_dfm_mx0[0])})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_qelse_conc_itm_33
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1[33:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2
      = ({1'b1 , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm[0])})
      + conv_u2s_34_35(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2[34:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva[32:0])
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_0})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_itm
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_mux_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2[0]),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_o000000
      = ~((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_lpi_2_dfm_34_1_mx0!=34'b0000000000000000000000000000000000)
      | (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_mux_nl));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl
      = conv_u2s_1_60(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_o000000)
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
      , operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_33_itm
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
      , operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_33_itm
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
      , operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_33_itm
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_33
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_33
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_33
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva[33])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp[33])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl[59:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13
      = readslicef_60_47_13((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_nl));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_lpi_2_dfm_34_1_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp,
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_sva_2[34:1]),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_47_tmp[33]);
  assign nl_quadInters_qnorm_rorig_run_acc_nl = conv_s2s_47_48(quadInters_qnorm_rorig_run_mul_1_cmp_4_z_oreg[46:0])
      + conv_s2s_47_48(quadInters_qnorm_rorig_run_mul_1_cmp_z_oreg[46:0]) + conv_s2s_47_48(quadInters_qnorm_rorig_run_mul_1_cmp_5_z_oreg[46:0]);
  assign quadInters_qnorm_rorig_run_acc_nl = nl_quadInters_qnorm_rorig_run_acc_nl[47:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1
      = conv_s2s_31_34(quads_crt_sva_1_376_112[183:153]) - (readslicef_48_34_14((quadInters_qnorm_rorig_run_acc_nl)));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_dividend_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      z_out_6[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_60_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_59_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_58_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_38_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_38_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_38_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_39_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_37_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1[32:0])
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_37_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_38_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_36_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva[32:0])
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_36_nl)
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_40_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_39_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_38_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_35_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      z_out_10[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1
      = ({(z_out_10[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[15])})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_12_cse
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_35_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1[34:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1
      = conv_u2s_1_34(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx0_33_32[1])
      + div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_64_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_64_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_64_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_65_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_63_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_63_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_63_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_64_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_62_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1
      = ({reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd_1
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_62_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_63_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33:0];
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1
      = ({(z_out_6[32:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_66_lpi_2_dfm_mx0[0])})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_qelse_conc_itm_33
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_68_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_66_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_65_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_64_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_63_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_44_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_44_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_44_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_45_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_43_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[32:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_43_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_43_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_44_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_42_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (z_out_7[33]));
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1
      = ({(z_out_7[32:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_42_lpi_2_dfm_mx0[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_42_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_43_lpi_2_dfm_mx0[33:1])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_46_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_45_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_44_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_43_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      z_out_7[33]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_42_lpi_2_dfm_mx0
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_24_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_49_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1[33:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[8])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_24_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_49_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_47_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      z_out_9[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1
      = ({(z_out_9[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[9])})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_13_cse
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_47_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_80_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1[33:0])
      , (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[28])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_80_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_7_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_3_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_81_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1[33:0])
      , (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[29])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_3_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_81_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_6_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_2_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_82_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1[33:0])
      , (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[30])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_2_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_82_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_5_sva_1[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_1_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_83_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[33:0])
      , (quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[31])}) + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_1_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_83_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_4_sva_1[34:0];
  assign for_nor_tmp = ~(for_stage_0 | for_stage_0_1 | for_stage_0_2 | for_stage_0_3
      | for_stage_0_4 | for_stage_0_5 | for_stage_0_6 | for_stage_0_7 | for_stage_0_8
      | for_stage_0_9);
  assign nl_quadInters_run_if_1_acc_nl = conv_s2u_34_35(ac_math_ac_abs_58_58_xabs_57_24_sva)
      + 35'b11111111111111111111111111111111111;
  assign quadInters_run_if_1_acc_nl = nl_quadInters_run_if_1_acc_nl[34:0];
  assign quadInters_run_if_1_acc_itm_34 = readslicef_35_1_34((quadInters_run_if_1_acc_nl));
  assign quadInters_run_mux_593_tmp_33 = MUX_s_1_2_2((quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56[1]),
      (quadInters_run_if_1_exs_mx1w0_1_0[1]), quadInters_run_if_1_acc_itm_34);
  assign and_dcpl_54 = (~(quadInters_run_land_lpi_2_dfm_st_7 | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6))
      & for_stage_0_8;
  assign or_69_cse = quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 | quadInters_run_land_lpi_2_dfm_8
      | quadInters_run_lor_lpi_2_dfm_1;
  assign and_dcpl_195 = for_stage_0_7 & (~ quadInters_run_land_lpi_2_dfm_st_6) &
      (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_5);
  assign or_dcpl_79 = (fsm_output[4:3]!=2'b00);
  assign and_dcpl_200 = ~((fsm_output[0]) | (fsm_output[6]));
  assign or_dcpl_91 = (fsm_output[0]) | (fsm_output[6]);
  assign or_dcpl_95 = operator_33_true_asn_1_itm_8 | (~ for_stage_0_9);
  assign and_dcpl_238 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2
      & for_stage_0_4 & (~(quadInters_run_land_lpi_2_dfm_st_3 | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2));
  assign or_tmp_328 = (quadInters_run_if_5_quadInters_run_if_5_or_2_tmp | or_69_cse)
      & for_stage_0_9 & (fsm_output[2]);
  assign or_tmp_480 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
      & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st
      & (fsm_output[3]);
  assign or_tmp_481 = div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st)
      & (fsm_output[3]);
  assign or_tmp_490 = (~ for_hitWorld_lpi_2_dfm_2) & for_stage_0_9 & (fsm_output[3]);
  assign or_tmp_529 = or_dcpl_91 | (fsm_output[1]);
  assign and_1128_cse = or_1462_cse | (fsm_output[3]);
  assign or_tmp_531 = and_1128_cse | ((quadInters_run_if_5_quadInters_run_if_5_or_2_tmp
      | or_69_cse | or_dcpl_95) & (fsm_output[2]));
  assign or_tmp_673 = ((operator_33_true_asn_1_itm_8 | (~ for_hitWorld_lpi_2_dfm_2)
      | (~ for_stage_0_9)) & (fsm_output[3])) | or_1462_cse | (fsm_output[2]);
  assign or_tmp_691 = and_dcpl_200 & (~ (fsm_output[1]));
  assign operator_33_true_asn_1_itm_9_mx0c2 = for_stage_0_9 & (fsm_output[5]);
  assign mult_run_mul_cmp_a = MUX1HOT_v_34_3_2((ray_temp_in_crt_sva[130:97]), (ray_temp_in_crt_sva[96:63]),
      (ray_temp_in_crt_sva[164:131]), {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[5])});
  assign mult_run_mul_cmp_b = {quadInters_run_t_trunc_mux_47_cse , quadInters_run_t_trunc_mux_48_cse
      , quadInters_run_t_trunc_mux_49_cse , quadInters_run_t_trunc_mux_50_cse , quadInters_run_t_trunc_mux_51_cse
      , quadInters_run_t_trunc_mux_52_cse , quadInters_run_t_trunc_mux_53_cse , quadInters_run_t_trunc_mux_54_cse
      , quadInters_run_t_trunc_mux_55_cse , quadInters_run_t_trunc_mux_56_cse , quadInters_run_t_trunc_mux_57_cse
      , quadInters_run_t_trunc_mux_58_cse , quadInters_run_t_trunc_mux_59_cse , quadInters_run_t_trunc_mux_60_cse
      , quadInters_run_t_trunc_mux_61_cse , quadInters_run_t_trunc_mux_62_cse , quadInters_run_t_trunc_mux_63_cse
      , quadInters_run_t_trunc_mux_64_cse , quadInters_run_t_trunc_mux_65_cse , quadInters_run_t_trunc_mux_66_cse
      , quadInters_run_t_trunc_mux_67_cse , quadInters_run_t_trunc_mux_68_cse , quadInters_run_t_trunc_mux_69_cse
      , quadInters_run_t_trunc_mux_70_cse , quadInters_run_t_trunc_mux_71_cse , quadInters_run_t_trunc_mux_72_cse
      , quadInters_run_t_trunc_mux_73_cse , quadInters_run_t_trunc_mux_74_cse , quadInters_run_t_trunc_mux_75_cse
      , quadInters_run_t_trunc_mux_76_cse , quadInters_run_t_trunc_mux_77_cse , quadInters_run_t_trunc_mux_78_cse
      , quadInters_run_t_trunc_mux_79_cse , quadInters_run_t_trunc_mux_80_cse , quadInters_run_t_trunc_mux_81_cse
      , quadInters_run_t_trunc_mux_82_cse , quadInters_run_t_trunc_mux_83_cse , quadInters_run_t_trunc_mux_84_cse
      , quadInters_run_t_trunc_mux_85_cse , quadInters_run_t_trunc_mux_86_cse , quadInters_run_t_trunc_mux_87_cse
      , quadInters_run_t_trunc_mux_88_cse , quadInters_run_t_trunc_mux_89_cse , quadInters_run_t_trunc_mux_90_cse
      , quadInters_run_t_trunc_mux_91_cse , quadInters_run_t_trunc_mux_92_cse , quadInters_run_t_trunc_mux_93_cse};
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_mux_10_itm
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      z_out_4[33]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_out_rsci_idat_0 <= 1'b0;
      closest_so_far_out_rsci_idat_1 <= 1'b0;
      closest_so_far_out_rsci_idat_2 <= 1'b0;
      closest_so_far_out_rsci_idat_3 <= 1'b0;
      closest_so_far_out_rsci_idat_4 <= 1'b0;
      closest_so_far_out_rsci_idat_5 <= 1'b0;
      closest_so_far_out_rsci_idat_6 <= 1'b0;
      closest_so_far_out_rsci_idat_7 <= 1'b0;
      closest_so_far_out_rsci_idat_8 <= 1'b0;
      closest_so_far_out_rsci_idat_9 <= 1'b0;
      closest_so_far_out_rsci_idat_10 <= 1'b0;
      closest_so_far_out_rsci_idat_11 <= 1'b0;
      closest_so_far_out_rsci_idat_12 <= 1'b0;
      closest_so_far_out_rsci_idat_13 <= 1'b0;
      closest_so_far_out_rsci_idat_14 <= 1'b0;
      closest_so_far_out_rsci_idat_15 <= 1'b0;
      closest_so_far_out_rsci_idat_16 <= 1'b0;
      closest_so_far_out_rsci_idat_17 <= 1'b0;
      closest_so_far_out_rsci_idat_18 <= 1'b0;
      closest_so_far_out_rsci_idat_19 <= 1'b0;
      closest_so_far_out_rsci_idat_20 <= 1'b0;
      closest_so_far_out_rsci_idat_21 <= 1'b0;
      closest_so_far_out_rsci_idat_22 <= 1'b0;
      closest_so_far_out_rsci_idat_23 <= 1'b0;
      closest_so_far_out_rsci_idat_24 <= 1'b0;
      closest_so_far_out_rsci_idat_25 <= 1'b0;
      closest_so_far_out_rsci_idat_26 <= 1'b0;
      closest_so_far_out_rsci_idat_27 <= 1'b0;
      closest_so_far_out_rsci_idat_28 <= 1'b0;
      closest_so_far_out_rsci_idat_29 <= 1'b0;
      closest_so_far_out_rsci_idat_30 <= 1'b0;
      closest_so_far_out_rsci_idat_31 <= 1'b0;
      closest_so_far_out_rsci_idat_32 <= 1'b0;
      closest_so_far_out_rsci_idat_33 <= 1'b0;
      closest_so_far_out_rsci_idat_34 <= 1'b0;
      closest_so_far_out_rsci_idat_35 <= 1'b0;
      closest_so_far_out_rsci_idat_36 <= 1'b0;
      closest_so_far_out_rsci_idat_37 <= 1'b0;
      closest_so_far_out_rsci_idat_38 <= 1'b0;
      closest_so_far_out_rsci_idat_39 <= 1'b0;
      closest_so_far_out_rsci_idat_40 <= 1'b0;
      closest_so_far_out_rsci_idat_41 <= 1'b0;
      closest_so_far_out_rsci_idat_42 <= 1'b0;
      closest_so_far_out_rsci_idat_43 <= 1'b0;
      closest_so_far_out_rsci_idat_44 <= 1'b0;
      closest_so_far_out_rsci_idat_45 <= 1'b0;
      closest_so_far_out_rsci_idat_46 <= 1'b0;
      rec_quad_out_rsci_idat_0 <= 1'b0;
      rec_quad_out_rsci_idat_20_1 <= 20'b00000000000000000000;
      rec_quad_out_rsci_idat_21 <= 1'b0;
      rec_quad_out_rsci_idat_41_22 <= 20'b00000000000000000000;
      rec_quad_out_rsci_idat_42 <= 1'b0;
      rec_quad_out_rsci_idat_62_43 <= 20'b00000000000000000000;
      rec_quad_out_rsci_idat_88_63 <= 26'b00000000000000000000000000;
      rec_quad_out_rsci_idat_114_89 <= 26'b00000000000000000000000000;
      rec_quad_out_rsci_idat_140_115 <= 26'b00000000000000000000000000;
      rec_quad_out_rsci_idat_141 <= 1'b0;
      rec_quad_out_rsci_idat_144_142 <= 3'b000;
      rec_quad_out_rsci_idat_171_145 <= 27'b000000000000000000000000000;
      rec_quad_out_rsci_idat_198_172 <= 27'b000000000000000000000000000;
      rec_quad_out_rsci_idat_225_199 <= 27'b000000000000000000000000000;
      quad_hit_anything_out_rsci_idat <= 1'b0;
    end
    else if ( closest_so_far_out_and_cse ) begin
      closest_so_far_out_rsci_idat_0 <= closest_so_far_sva_dfm_3_0;
      closest_so_far_out_rsci_idat_1 <= closest_so_far_sva_dfm_3_1;
      closest_so_far_out_rsci_idat_2 <= closest_so_far_sva_dfm_3_2;
      closest_so_far_out_rsci_idat_3 <= closest_so_far_sva_dfm_3_3;
      closest_so_far_out_rsci_idat_4 <= closest_so_far_sva_dfm_3_4;
      closest_so_far_out_rsci_idat_5 <= closest_so_far_sva_dfm_3_5;
      closest_so_far_out_rsci_idat_6 <= closest_so_far_sva_dfm_3_6;
      closest_so_far_out_rsci_idat_7 <= closest_so_far_sva_dfm_3_7;
      closest_so_far_out_rsci_idat_8 <= closest_so_far_sva_dfm_3_8;
      closest_so_far_out_rsci_idat_9 <= closest_so_far_sva_dfm_3_9;
      closest_so_far_out_rsci_idat_10 <= closest_so_far_sva_dfm_3_10;
      closest_so_far_out_rsci_idat_11 <= closest_so_far_sva_dfm_3_11;
      closest_so_far_out_rsci_idat_12 <= closest_so_far_sva_dfm_3_12;
      closest_so_far_out_rsci_idat_13 <= closest_so_far_sva_dfm_3_13;
      closest_so_far_out_rsci_idat_14 <= closest_so_far_sva_dfm_3_14;
      closest_so_far_out_rsci_idat_15 <= closest_so_far_sva_dfm_3_15;
      closest_so_far_out_rsci_idat_16 <= closest_so_far_sva_dfm_3_16;
      closest_so_far_out_rsci_idat_17 <= closest_so_far_sva_dfm_3_17;
      closest_so_far_out_rsci_idat_18 <= closest_so_far_sva_dfm_3_18;
      closest_so_far_out_rsci_idat_19 <= closest_so_far_sva_dfm_3_19;
      closest_so_far_out_rsci_idat_20 <= closest_so_far_sva_dfm_3_20;
      closest_so_far_out_rsci_idat_21 <= closest_so_far_sva_dfm_3_21;
      closest_so_far_out_rsci_idat_22 <= closest_so_far_sva_dfm_3_22;
      closest_so_far_out_rsci_idat_23 <= closest_so_far_sva_dfm_3_23;
      closest_so_far_out_rsci_idat_24 <= closest_so_far_sva_dfm_3_24;
      closest_so_far_out_rsci_idat_25 <= closest_so_far_sva_dfm_3_25;
      closest_so_far_out_rsci_idat_26 <= closest_so_far_sva_dfm_3_26;
      closest_so_far_out_rsci_idat_27 <= closest_so_far_sva_dfm_3_27;
      closest_so_far_out_rsci_idat_28 <= closest_so_far_sva_dfm_3_28;
      closest_so_far_out_rsci_idat_29 <= closest_so_far_sva_dfm_3_29;
      closest_so_far_out_rsci_idat_30 <= closest_so_far_sva_dfm_3_30;
      closest_so_far_out_rsci_idat_31 <= closest_so_far_sva_dfm_3_31;
      closest_so_far_out_rsci_idat_32 <= closest_so_far_sva_dfm_3_32;
      closest_so_far_out_rsci_idat_33 <= closest_so_far_sva_dfm_3_33;
      closest_so_far_out_rsci_idat_34 <= closest_so_far_sva_dfm_3_34;
      closest_so_far_out_rsci_idat_35 <= closest_so_far_sva_dfm_3_35;
      closest_so_far_out_rsci_idat_36 <= closest_so_far_sva_dfm_3_36;
      closest_so_far_out_rsci_idat_37 <= closest_so_far_sva_dfm_3_37;
      closest_so_far_out_rsci_idat_38 <= closest_so_far_sva_dfm_3_38;
      closest_so_far_out_rsci_idat_39 <= closest_so_far_sva_dfm_3_39;
      closest_so_far_out_rsci_idat_40 <= closest_so_far_sva_dfm_3_40;
      closest_so_far_out_rsci_idat_41 <= closest_so_far_sva_dfm_3_41;
      closest_so_far_out_rsci_idat_42 <= closest_so_far_sva_dfm_3_42;
      closest_so_far_out_rsci_idat_43 <= closest_so_far_sva_dfm_3_43;
      closest_so_far_out_rsci_idat_44 <= closest_so_far_sva_dfm_3_44;
      closest_so_far_out_rsci_idat_45 <= closest_so_far_sva_dfm_3_45;
      closest_so_far_out_rsci_idat_46 <= closest_so_far_sva_dfm_3_46;
      rec_quad_out_rsci_idat_0 <= rec_quad_hit_loc_x_0_sva_dfm;
      rec_quad_out_rsci_idat_20_1 <= reg_ac_math_ac_abs_21_21_1_xabs_xor_ftd_1;
      rec_quad_out_rsci_idat_21 <= rec_quad_hit_loc_y_0_sva_dfm;
      rec_quad_out_rsci_idat_41_22 <= reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1;
      rec_quad_out_rsci_idat_42 <= rec_quad_hit_loc_z_0_sva_dfm;
      rec_quad_out_rsci_idat_62_43 <= reg_ac_math_ac_abs_21_21_xabs_xor_ftd_1;
      rec_quad_out_rsci_idat_88_63 <= rec_quad_normal_x_sva_dfm;
      rec_quad_out_rsci_idat_114_89 <= rec_quad_normal_y_sva_dfm;
      rec_quad_out_rsci_idat_140_115 <= rec_quad_normal_z_sva_dfm;
      rec_quad_out_rsci_idat_141 <= operator_33_true_asn_1_itm_9;
      rec_quad_out_rsci_idat_144_142 <= quads_crt_sva_8_110_108;
      rec_quad_out_rsci_idat_171_145 <= rec_quad_color_r_sva_dfm;
      rec_quad_out_rsci_idat_198_172 <= rec_quad_color_g_sva_dfm;
      rec_quad_out_rsci_idat_225_199 <= rec_quad_color_b_sva_dfm;
      quad_hit_anything_out_rsci_idat <= quad_hit_anything_sva_dfm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ensig_cgo <= 1'b0;
      reg_closest_so_far_out_rsci_ivld_hit_psct_cse <= 1'b0;
      reg_quad_max_in_rsci_irdy_hit_psct_cse <= 1'b0;
      reg_quads_rsci_irdy_hit_psct_cse <= 1'b0;
      quadInters_denom_dot_run_mul_1_cmp_b <= 34'b0000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_1_cmp_a <= 26'b00000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_1_b <= 34'b0000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_1_a <= 26'b00000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_b <= 34'b0000000000000000000000000000000000;
      quadInters_denom_dot_run_mul_2_cmp_a <= 26'b00000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_5_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_5_a <= 25'b0000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_4_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_4_a <= 25'b0000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_3_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_3_a <= 25'b0000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_2_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_2_a <= 25'b0000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_1_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_1_a <= 25'b0000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_b <= 56'b00000000000000000000000000000000000000000000000000000000;
      quadInters_qnorm_rorig_run_mul_1_cmp_a <= 25'b0000000000000000000000000;
      closest_so_far_sva_46 <= 1'b0;
      closest_so_far_sva_0 <= 1'b0;
      closest_so_far_sva_45 <= 1'b0;
      closest_so_far_sva_1 <= 1'b0;
      closest_so_far_sva_44 <= 1'b0;
      closest_so_far_sva_2 <= 1'b0;
      closest_so_far_sva_43 <= 1'b0;
      closest_so_far_sva_3 <= 1'b0;
      closest_so_far_sva_42 <= 1'b0;
      closest_so_far_sva_4 <= 1'b0;
      closest_so_far_sva_41 <= 1'b0;
      closest_so_far_sva_5 <= 1'b0;
      closest_so_far_sva_40 <= 1'b0;
      closest_so_far_sva_6 <= 1'b0;
      closest_so_far_sva_39 <= 1'b0;
      closest_so_far_sva_7 <= 1'b0;
      closest_so_far_sva_38 <= 1'b0;
      closest_so_far_sva_8 <= 1'b0;
      closest_so_far_sva_37 <= 1'b0;
      closest_so_far_sva_9 <= 1'b0;
      closest_so_far_sva_36 <= 1'b0;
      closest_so_far_sva_10 <= 1'b0;
      closest_so_far_sva_35 <= 1'b0;
      closest_so_far_sva_11 <= 1'b0;
      closest_so_far_sva_34 <= 1'b0;
      closest_so_far_sva_12 <= 1'b0;
      closest_so_far_sva_33 <= 1'b0;
      closest_so_far_sva_13 <= 1'b0;
      closest_so_far_sva_32 <= 1'b0;
      closest_so_far_sva_14 <= 1'b0;
      closest_so_far_sva_31 <= 1'b0;
      closest_so_far_sva_15 <= 1'b0;
      closest_so_far_sva_30 <= 1'b0;
      closest_so_far_sva_16 <= 1'b0;
      closest_so_far_sva_29 <= 1'b0;
      closest_so_far_sva_17 <= 1'b0;
      closest_so_far_sva_28 <= 1'b0;
      closest_so_far_sva_18 <= 1'b0;
      closest_so_far_sva_27 <= 1'b0;
      closest_so_far_sva_19 <= 1'b0;
      closest_so_far_sva_26 <= 1'b0;
      closest_so_far_sva_20 <= 1'b0;
      closest_so_far_sva_25 <= 1'b0;
      closest_so_far_sva_21 <= 1'b0;
      closest_so_far_sva_24 <= 1'b0;
      closest_so_far_sva_22 <= 1'b0;
      closest_so_far_sva_23 <= 1'b0;
      rec_quad_hit_loc_z_0_sva <= 1'b0;
      rec_quad_hit_loc_y_0_sva <= 1'b0;
      rec_quad_hit_loc_x_0_sva <= 1'b0;
      ray_temp_in_crt_sva <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_8_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quad_hit_anything_sva <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_46 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_45 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_44 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_43 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_42 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_41 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_40 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_39 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_38 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_37 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_36 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_35 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_34 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_33 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_32 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_31 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_30 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_29 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_28 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_27 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_26 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_25 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_24 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_23 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_22 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_21 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_20 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_19 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_18 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_17 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_16 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_15 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_14 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_13 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_12 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_11 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_10 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_9 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_8 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_7 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_6 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_5 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_4 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_3 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_2 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_1 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_1_0 <= 1'b0;
      for_stage_0 <= 1'b0;
      rec_quad_front_face_sva <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_32_0
          <= 33'b000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22
          <= 5'b00000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_33_itm
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva
          <= 35'b00000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
          <= 1'b0;
      reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg <= 2'b00;
      reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg <= 2'b00;
      reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg <= 2'b00;
      mult_run_asn_1_itm_74_43 <= 32'b00000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_32_0
          <= 33'b000000000000000000000000000000000;
      ac_math_ac_abs_58_58_xabs_57_24_sva <= 34'b0000000000000000000000000000000000;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_1_cse
          <= 33'b000000000000000000000000000000000;
      quadInters_at_run_mult_result_x_74_30_sva_12_0 <= 13'b0000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_0
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_32_0
          <= 33'b000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva
          <= 34'b0000000000000000000000000000000000;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd
          <= 33'b000000000000000000000000000000000;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd_1
          <= 33'b000000000000000000000000000000000;
    end
    else if ( hit_wen ) begin
      ensig_cgo <= ensig_cgo_mx0;
      reg_closest_so_far_out_rsci_ivld_hit_psct_cse <= for_nor_tmp & (fsm_output[5]);
      reg_quad_max_in_rsci_irdy_hit_psct_cse <= ~ and_dcpl_200;
      reg_quads_rsci_irdy_hit_psct_cse <= (for_stage_0 & (fsm_output[5])) | (fsm_output[1]);
      quadInters_denom_dot_run_mul_1_cmp_b <= MUX1HOT_v_34_3_2((ray_temp_in_crt_sva[130:97]),
          (ray_temp_in_crt_sva[164:131]), (ray_temp_in_crt_sva[96:63]), {or_cse ,
          (fsm_output[4]) , (fsm_output[5])});
      quadInters_denom_dot_run_mul_1_cmp_a <= MUX1HOT_v_26_4_2((quads_rsci_idat_mxwt[163:138]),
          (quads_crt_sva_8_189_112[51:26]), (quads_crt_sva_8_189_112[77:52]), (quads_crt_sva_8_189_112[25:0]),
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
      quadInters_denom_dot_run_mul_2_cmp_1_b <= ray_temp_in_crt_sva[96:63];
      quadInters_denom_dot_run_mul_2_cmp_1_a <= quads_rsci_idat_mxwt[137:112];
      quadInters_denom_dot_run_mul_2_cmp_b <= ray_temp_in_crt_sva[164:131];
      quadInters_denom_dot_run_mul_2_cmp_a <= quads_rsci_idat_mxwt[189:164];
      quadInters_qnorm_rorig_run_mul_1_cmp_5_b <= MUX_v_56_2_2((signext_56_26(quads_crt_sva_1_376_112[77:52])),
          (readslicef_57_56_1((quadInters_cross_u_run_acc_nl))), fsm_output[4]);
      quadInters_qnorm_rorig_run_mul_1_cmp_5_a <= MUX_v_25_2_2((signext_25_21(ray_temp_in_crt_sva[62:42])),
          (quads_crt_sva_7_264_112[102:78]), fsm_output[4]);
      quadInters_qnorm_rorig_run_mul_1_cmp_4_b <= MUX_v_56_2_2((signext_56_26(quads_crt_sva_1_376_112[25:0])),
          (readslicef_57_56_1((quadInters_cross_u_run_acc_2_nl))), fsm_output[4]);
      quadInters_qnorm_rorig_run_mul_1_cmp_4_a <= MUX_v_25_2_2((signext_25_21(ray_temp_in_crt_sva[20:0])),
          (quads_crt_sva_7_264_112[152:128]), fsm_output[4]);
      quadInters_qnorm_rorig_run_mul_1_cmp_3_b <= readslicef_57_56_1((quadInters_cross_v_run_acc_2_nl));
      quadInters_qnorm_rorig_run_mul_1_cmp_3_a <= quads_crt_sva_7_264_112[152:128];
      quadInters_qnorm_rorig_run_mul_1_cmp_2_b <= readslicef_57_56_1((quadInters_cross_v_run_acc_nl));
      quadInters_qnorm_rorig_run_mul_1_cmp_2_a <= quads_crt_sva_7_264_112[102:78];
      quadInters_qnorm_rorig_run_mul_1_cmp_1_b <= readslicef_57_56_1((quadInters_cross_u_run_acc_1_nl));
      quadInters_qnorm_rorig_run_mul_1_cmp_1_a <= quads_crt_sva_7_264_112[127:103];
      quadInters_qnorm_rorig_run_mul_1_cmp_b <= MUX_v_56_2_2((signext_56_26(quads_crt_sva_1_376_112[51:26])),
          (z_out[56:1]), fsm_output[4]);
      quadInters_qnorm_rorig_run_mul_1_cmp_a <= MUX_v_25_2_2((signext_25_21(ray_temp_in_crt_sva[41:21])),
          (quads_crt_sva_7_264_112[127:103]), fsm_output[4]);
      closest_so_far_sva_46 <= (quad_hit_anything_mux_48_nl) & (~ or_tmp_529);
      closest_so_far_sva_0 <= (quad_hit_anything_mux_47_nl) & (~ or_tmp_529);
      closest_so_far_sva_45 <= (quad_hit_anything_mux_46_nl) & (~ or_tmp_529);
      closest_so_far_sva_1 <= (quad_hit_anything_mux_45_nl) & (~ or_tmp_529);
      closest_so_far_sva_44 <= (quad_hit_anything_mux_44_nl) & (~ or_tmp_529);
      closest_so_far_sva_2 <= (quad_hit_anything_mux_43_nl) & (~ or_tmp_529);
      closest_so_far_sva_43 <= (quad_hit_anything_mux_42_nl) & (~ or_tmp_529);
      closest_so_far_sva_3 <= (quad_hit_anything_mux_41_nl) & (~ or_tmp_529);
      closest_so_far_sva_42 <= (quad_hit_anything_mux_40_nl) & (~ or_tmp_529);
      closest_so_far_sva_4 <= (quad_hit_anything_mux_39_nl) & (~ or_tmp_529);
      closest_so_far_sva_41 <= (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_4_nl)
          | or_tmp_529;
      closest_so_far_sva_5 <= (quad_hit_anything_mux_38_nl) & (~ or_tmp_529);
      closest_so_far_sva_40 <= (quad_hit_anything_mux_37_nl) & (~ or_tmp_529);
      closest_so_far_sva_6 <= (quad_hit_anything_mux_36_nl) & (~ or_tmp_529);
      closest_so_far_sva_39 <= (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_3_nl)
          | or_tmp_529;
      closest_so_far_sva_7 <= (quad_hit_anything_mux_35_nl) & (~ or_tmp_529);
      closest_so_far_sva_38 <= (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_2_nl)
          | or_tmp_529;
      closest_so_far_sva_8 <= (quad_hit_anything_mux_34_nl) & (~ or_tmp_529);
      closest_so_far_sva_37 <= (quad_hit_anything_mux_33_nl) & (~ or_tmp_529);
      closest_so_far_sva_9 <= (quad_hit_anything_mux_32_nl) & (~ or_tmp_529);
      closest_so_far_sva_36 <= (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_1_nl)
          | or_tmp_529;
      closest_so_far_sva_10 <= (quad_hit_anything_mux_31_nl) & (~ or_tmp_529);
      closest_so_far_sva_35 <= (quad_hit_anything_mux_30_nl) & (~ or_tmp_529);
      closest_so_far_sva_11 <= (quad_hit_anything_mux_29_nl) & (~ or_tmp_529);
      closest_so_far_sva_34 <= (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_nl)
          | or_tmp_529;
      closest_so_far_sva_12 <= (quad_hit_anything_mux_28_nl) & (~ or_tmp_529);
      closest_so_far_sva_33 <= (quad_hit_anything_mux_27_nl) & (~ or_tmp_529);
      closest_so_far_sva_13 <= (quad_hit_anything_mux_26_nl) & (~ or_tmp_529);
      closest_so_far_sva_32 <= (quad_hit_anything_mux_25_nl) & (~ or_tmp_529);
      closest_so_far_sva_14 <= (quad_hit_anything_mux_24_nl) & (~ or_tmp_529);
      closest_so_far_sva_31 <= (quad_hit_anything_mux_23_nl) & (~ or_tmp_529);
      closest_so_far_sva_15 <= (quad_hit_anything_mux_22_nl) & (~ or_tmp_529);
      closest_so_far_sva_30 <= (quad_hit_anything_mux_21_nl) & (~ or_tmp_529);
      closest_so_far_sva_16 <= (quad_hit_anything_mux_20_nl) & (~ or_tmp_529);
      closest_so_far_sva_29 <= (quad_hit_anything_mux_19_nl) & (~ or_tmp_529);
      closest_so_far_sva_17 <= (quad_hit_anything_mux_18_nl) & (~ or_tmp_529);
      closest_so_far_sva_28 <= (quad_hit_anything_mux_17_nl) & (~ or_tmp_529);
      closest_so_far_sva_18 <= (quad_hit_anything_mux_16_nl) & (~ or_tmp_529);
      closest_so_far_sva_27 <= (quad_hit_anything_mux_15_nl) & (~ or_tmp_529);
      closest_so_far_sva_19 <= (quad_hit_anything_mux_14_nl) & (~ or_tmp_529);
      closest_so_far_sva_26 <= (quad_hit_anything_mux_13_nl) & (~ or_tmp_529);
      closest_so_far_sva_20 <= (quad_hit_anything_mux_12_nl) & (~ or_tmp_529);
      closest_so_far_sva_25 <= (quad_hit_anything_mux_11_nl) & (~ or_tmp_529);
      closest_so_far_sva_21 <= (quad_hit_anything_mux_10_nl) & (~ or_tmp_529);
      closest_so_far_sva_24 <= (quad_hit_anything_mux_9_nl) & (~ or_tmp_529);
      closest_so_far_sva_22 <= (quad_hit_anything_mux_8_nl) & (~ or_tmp_529);
      closest_so_far_sva_23 <= (quad_hit_anything_mux_7_nl) & (~ or_tmp_529);
      rec_quad_hit_loc_z_0_sva <= (quad_hit_anything_mux_6_nl) & (~ or_tmp_529);
      rec_quad_hit_loc_y_0_sva <= (quad_hit_anything_mux_5_nl) & (~ or_tmp_529);
      rec_quad_hit_loc_x_0_sva <= (quad_hit_anything_mux_4_nl) & (~ or_tmp_529);
      ray_temp_in_crt_sva <= MUX_v_166_2_2(ray_temp_in_rsci_idat_mxwt, ray_temp_in_crt_sva,
          or_tmp_691);
      quads_crt_sva_8_376_296 <= quads_crt_sva_7_376_296;
      quad_hit_anything_sva <= (quad_hit_anything_mux_nl) & (~ or_tmp_529);
      quadInters_run_t_trunc_lpi_2_dfm_1_46 <= quadInters_run_t_trunc_mux_47_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_45 <= quadInters_run_t_trunc_mux_48_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_44 <= quadInters_run_t_trunc_mux_49_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_43 <= quadInters_run_t_trunc_mux_50_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_42 <= quadInters_run_t_trunc_mux_51_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_41 <= quadInters_run_t_trunc_mux_52_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_40 <= quadInters_run_t_trunc_mux_53_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_39 <= quadInters_run_t_trunc_mux_54_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_38 <= quadInters_run_t_trunc_mux_55_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_37 <= quadInters_run_t_trunc_mux_56_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_36 <= quadInters_run_t_trunc_mux_57_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_35 <= quadInters_run_t_trunc_mux_58_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_34 <= quadInters_run_t_trunc_mux_59_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_33 <= quadInters_run_t_trunc_mux_60_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_32 <= quadInters_run_t_trunc_mux_61_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_31 <= quadInters_run_t_trunc_mux_62_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_30 <= quadInters_run_t_trunc_mux_63_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_29 <= quadInters_run_t_trunc_mux_64_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_28 <= quadInters_run_t_trunc_mux_65_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_27 <= quadInters_run_t_trunc_mux_66_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_26 <= quadInters_run_t_trunc_mux_67_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_25 <= quadInters_run_t_trunc_mux_68_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_24 <= quadInters_run_t_trunc_mux_69_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_23 <= quadInters_run_t_trunc_mux_70_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_22 <= quadInters_run_t_trunc_mux_71_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_21 <= quadInters_run_t_trunc_mux_72_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_20 <= quadInters_run_t_trunc_mux_73_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_19 <= quadInters_run_t_trunc_mux_74_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_18 <= quadInters_run_t_trunc_mux_75_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_17 <= quadInters_run_t_trunc_mux_76_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_16 <= quadInters_run_t_trunc_mux_77_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_15 <= quadInters_run_t_trunc_mux_78_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_14 <= quadInters_run_t_trunc_mux_79_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_13 <= quadInters_run_t_trunc_mux_80_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_12 <= quadInters_run_t_trunc_mux_81_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_11 <= quadInters_run_t_trunc_mux_82_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_10 <= quadInters_run_t_trunc_mux_83_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_9 <= quadInters_run_t_trunc_mux_84_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_8 <= quadInters_run_t_trunc_mux_85_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_7 <= quadInters_run_t_trunc_mux_86_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_6 <= quadInters_run_t_trunc_mux_87_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_5 <= quadInters_run_t_trunc_mux_88_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_4 <= quadInters_run_t_trunc_mux_89_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_3 <= quadInters_run_t_trunc_mux_90_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_2 <= quadInters_run_t_trunc_mux_91_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_1 <= quadInters_run_t_trunc_mux_92_cse;
      quadInters_run_t_trunc_lpi_2_dfm_1_0 <= quadInters_run_t_trunc_mux_93_cse;
      for_stage_0 <= (for_stage_0 & (~(or_dcpl_91 | (or_343_cse & for_stage_0_1 &
          (fsm_output[2]))))) | (fsm_output[1]);
      rec_quad_front_face_sva <= (quad_hit_anything_mux_3_nl) & (~ or_tmp_529);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[0]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[1]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[10]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[11]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_3,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[12]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[13]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[14]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[15]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[16]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[17]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[18]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[19]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2
          <= MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_2,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[2]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1,
          {or_cse , operator_35_true_and_57_cse , operator_35_true_and_58_cse , (fsm_output[5])});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_32_0
          <= z_out_4[32:0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22
          <= quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[26:22];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_33_itm
          <= MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva
          <= MUX_v_35_2_2(z_out_3, z_out_8, div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_m1c);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs
          <= (quad_hit_anything_mux1h_58_nl) & (~ or_tmp_529);
      reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg <= quadInters_sub_run_mux_rgt[22:21];
      reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg <= quadInters_sub_run_mux_1_rgt[22:21];
      reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg <= quadInters_sub_run_mux_2_rgt[22:21];
      mult_run_asn_1_itm_74_43 <= mult_run_mul_cmp_z_oreg[44:13];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_32_0
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt[32:0];
      ac_math_ac_abs_58_58_xabs_57_24_sva <= MUX_v_34_2_2(ac_math_ac_abs_58_58_xabs_acc_itm_57_24,
          ({33'b000000000000000000000000000000000 , (ac_math_ac_abs_58_58_xabs_57_24_sva_mx1[0])}),
          fsm_output[3]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_1_cse
          <= z_out_2[32:0];
      quadInters_at_run_mult_result_x_74_30_sva_12_0 <= mult_run_mul_cmp_z_oreg[12:0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_nl),
          (operator_35_true_mux_172_nl), fsm_output[4]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_45_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_0
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_78_lpi_2_dfm_mx0[0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_44_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_43_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_32_0
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1[32:0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva
          <= MUX_v_34_2_2(z_out_4, div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1,
          fsm_output[4]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_mux_10_itm[33:1];
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1
          <= MUX1HOT_s_1_4_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx1[0]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx2[0]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx3[0]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_mux_10_itm[0]),
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_ftd_1
          <= MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_74_lpi_2_dfm_mx0[0]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_mux_10_itm[0]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_mx2[0]),
          {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd_1
          <= z_out_3[32:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      closest_so_far_sva_dfm_3_46 <= 1'b0;
      closest_so_far_sva_dfm_3_0 <= 1'b0;
      closest_so_far_sva_dfm_3_45 <= 1'b0;
      closest_so_far_sva_dfm_3_1 <= 1'b0;
      closest_so_far_sva_dfm_3_44 <= 1'b0;
      closest_so_far_sva_dfm_3_2 <= 1'b0;
      closest_so_far_sva_dfm_3_43 <= 1'b0;
      closest_so_far_sva_dfm_3_3 <= 1'b0;
      closest_so_far_sva_dfm_3_42 <= 1'b0;
      closest_so_far_sva_dfm_3_4 <= 1'b0;
      closest_so_far_sva_dfm_3_41 <= 1'b0;
      closest_so_far_sva_dfm_3_5 <= 1'b0;
      closest_so_far_sva_dfm_3_40 <= 1'b0;
      closest_so_far_sva_dfm_3_6 <= 1'b0;
      closest_so_far_sva_dfm_3_39 <= 1'b0;
      closest_so_far_sva_dfm_3_7 <= 1'b0;
      closest_so_far_sva_dfm_3_38 <= 1'b0;
      closest_so_far_sva_dfm_3_8 <= 1'b0;
      closest_so_far_sva_dfm_3_37 <= 1'b0;
      closest_so_far_sva_dfm_3_9 <= 1'b0;
      closest_so_far_sva_dfm_3_36 <= 1'b0;
      closest_so_far_sva_dfm_3_10 <= 1'b0;
      closest_so_far_sva_dfm_3_35 <= 1'b0;
      closest_so_far_sva_dfm_3_11 <= 1'b0;
      closest_so_far_sva_dfm_3_34 <= 1'b0;
      closest_so_far_sva_dfm_3_12 <= 1'b0;
      closest_so_far_sva_dfm_3_33 <= 1'b0;
      closest_so_far_sva_dfm_3_13 <= 1'b0;
      closest_so_far_sva_dfm_3_32 <= 1'b0;
      closest_so_far_sva_dfm_3_14 <= 1'b0;
      closest_so_far_sva_dfm_3_31 <= 1'b0;
      closest_so_far_sva_dfm_3_15 <= 1'b0;
      closest_so_far_sva_dfm_3_30 <= 1'b0;
      closest_so_far_sva_dfm_3_16 <= 1'b0;
      closest_so_far_sva_dfm_3_29 <= 1'b0;
      closest_so_far_sva_dfm_3_17 <= 1'b0;
      closest_so_far_sva_dfm_3_28 <= 1'b0;
      closest_so_far_sva_dfm_3_18 <= 1'b0;
      closest_so_far_sva_dfm_3_27 <= 1'b0;
      closest_so_far_sva_dfm_3_19 <= 1'b0;
      closest_so_far_sva_dfm_3_26 <= 1'b0;
      closest_so_far_sva_dfm_3_20 <= 1'b0;
      closest_so_far_sva_dfm_3_25 <= 1'b0;
      closest_so_far_sva_dfm_3_21 <= 1'b0;
      closest_so_far_sva_dfm_3_24 <= 1'b0;
      closest_so_far_sva_dfm_3_22 <= 1'b0;
      closest_so_far_sva_dfm_3_23 <= 1'b0;
    end
    else if ( closest_so_far_and_47_cse ) begin
      closest_so_far_sva_dfm_3_46 <= MUX_s_1_2_2(closest_so_far_sva_46, quadInters_run_t_trunc_lpi_2_dfm_2_46,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_0 <= MUX_s_1_2_2(closest_so_far_sva_0, quadInters_run_t_trunc_lpi_2_dfm_2_0,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_45 <= MUX_s_1_2_2(closest_so_far_sva_45, quadInters_run_t_trunc_lpi_2_dfm_2_45,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_1 <= MUX_s_1_2_2(closest_so_far_sva_1, quadInters_run_t_trunc_lpi_2_dfm_2_1,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_44 <= MUX_s_1_2_2(closest_so_far_sva_44, quadInters_run_t_trunc_lpi_2_dfm_2_44,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_2 <= MUX_s_1_2_2(closest_so_far_sva_2, quadInters_run_t_trunc_lpi_2_dfm_2_2,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_43 <= MUX_s_1_2_2(closest_so_far_sva_43, quadInters_run_t_trunc_lpi_2_dfm_2_43,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_3 <= MUX_s_1_2_2(closest_so_far_sva_3, quadInters_run_t_trunc_lpi_2_dfm_2_3,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_42 <= MUX_s_1_2_2(closest_so_far_sva_42, quadInters_run_t_trunc_lpi_2_dfm_2_42,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_4 <= MUX_s_1_2_2(closest_so_far_sva_4, quadInters_run_t_trunc_lpi_2_dfm_2_4,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_41 <= MUX_s_1_2_2(closest_so_far_sva_41, quadInters_run_t_trunc_lpi_2_dfm_2_41,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_5 <= MUX_s_1_2_2(closest_so_far_sva_5, quadInters_run_t_trunc_lpi_2_dfm_2_5,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_40 <= MUX_s_1_2_2(closest_so_far_sva_40, quadInters_run_t_trunc_lpi_2_dfm_2_40,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_6 <= MUX_s_1_2_2(closest_so_far_sva_6, quadInters_run_t_trunc_lpi_2_dfm_2_6,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_39 <= MUX_s_1_2_2(closest_so_far_sva_39, quadInters_run_t_trunc_lpi_2_dfm_2_39,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_7 <= MUX_s_1_2_2(closest_so_far_sva_7, quadInters_run_t_trunc_lpi_2_dfm_2_7,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_38 <= MUX_s_1_2_2(closest_so_far_sva_38, quadInters_run_t_trunc_lpi_2_dfm_2_38,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_8 <= MUX_s_1_2_2(closest_so_far_sva_8, quadInters_run_t_trunc_lpi_2_dfm_2_8,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_37 <= MUX_s_1_2_2(closest_so_far_sva_37, quadInters_run_t_trunc_lpi_2_dfm_2_37,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_9 <= MUX_s_1_2_2(closest_so_far_sva_9, quadInters_run_t_trunc_lpi_2_dfm_2_9,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_36 <= MUX_s_1_2_2(closest_so_far_sva_36, quadInters_run_t_trunc_lpi_2_dfm_2_36,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_10 <= MUX_s_1_2_2(closest_so_far_sva_10, quadInters_run_t_trunc_lpi_2_dfm_2_10,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_35 <= MUX_s_1_2_2(closest_so_far_sva_35, quadInters_run_t_trunc_lpi_2_dfm_2_35,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_11 <= MUX_s_1_2_2(closest_so_far_sva_11, quadInters_run_t_trunc_lpi_2_dfm_2_11,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_34 <= MUX_s_1_2_2(closest_so_far_sva_34, quadInters_run_t_trunc_lpi_2_dfm_2_34,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_12 <= MUX_s_1_2_2(closest_so_far_sva_12, quadInters_run_t_trunc_lpi_2_dfm_2_12,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_33 <= MUX_s_1_2_2(closest_so_far_sva_33, quadInters_run_t_trunc_lpi_2_dfm_2_33,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_13 <= MUX_s_1_2_2(closest_so_far_sva_13, quadInters_run_t_trunc_lpi_2_dfm_2_13,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_32 <= MUX_s_1_2_2(closest_so_far_sva_32, quadInters_run_t_trunc_lpi_2_dfm_2_32,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_14 <= MUX_s_1_2_2(closest_so_far_sva_14, quadInters_run_t_trunc_lpi_2_dfm_2_14,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_31 <= MUX_s_1_2_2(closest_so_far_sva_31, quadInters_run_t_trunc_lpi_2_dfm_2_31,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_15 <= MUX_s_1_2_2(closest_so_far_sva_15, quadInters_run_t_trunc_lpi_2_dfm_2_15,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_30 <= MUX_s_1_2_2(closest_so_far_sva_30, quadInters_run_t_trunc_lpi_2_dfm_2_30,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_16 <= MUX_s_1_2_2(closest_so_far_sva_16, quadInters_run_t_trunc_lpi_2_dfm_2_16,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_29 <= MUX_s_1_2_2(closest_so_far_sva_29, quadInters_run_t_trunc_lpi_2_dfm_2_29,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_17 <= MUX_s_1_2_2(closest_so_far_sva_17, quadInters_run_t_trunc_lpi_2_dfm_2_17,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_28 <= MUX_s_1_2_2(closest_so_far_sva_28, quadInters_run_t_trunc_lpi_2_dfm_2_28,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_18 <= MUX_s_1_2_2(closest_so_far_sva_18, quadInters_run_t_trunc_lpi_2_dfm_2_18,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_27 <= MUX_s_1_2_2(closest_so_far_sva_27, quadInters_run_t_trunc_lpi_2_dfm_2_27,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_19 <= MUX_s_1_2_2(closest_so_far_sva_19, quadInters_run_t_trunc_lpi_2_dfm_2_19,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_26 <= MUX_s_1_2_2(closest_so_far_sva_26, quadInters_run_t_trunc_lpi_2_dfm_2_26,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_20 <= MUX_s_1_2_2(closest_so_far_sva_20, quadInters_run_t_trunc_lpi_2_dfm_2_20,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_25 <= MUX_s_1_2_2(closest_so_far_sva_25, quadInters_run_t_trunc_lpi_2_dfm_2_25,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_21 <= MUX_s_1_2_2(closest_so_far_sva_21, quadInters_run_t_trunc_lpi_2_dfm_2_21,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_24 <= MUX_s_1_2_2(closest_so_far_sva_24, quadInters_run_t_trunc_lpi_2_dfm_2_24,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_22 <= MUX_s_1_2_2(closest_so_far_sva_22, quadInters_run_t_trunc_lpi_2_dfm_2_22,
          fsm_output[5]);
      closest_so_far_sva_dfm_3_23 <= MUX_s_1_2_2(closest_so_far_sva_23, quadInters_run_t_trunc_lpi_2_dfm_2_23,
          fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_color_b_sva_dfm <= 27'b000000000000000000000000000;
      rec_quad_color_g_sva_dfm <= 27'b000000000000000000000000000;
      rec_quad_color_r_sva_dfm <= 27'b000000000000000000000000000;
    end
    else if ( rec_quad_color_b_and_cse ) begin
      rec_quad_color_b_sva_dfm <= MUX_v_27_2_2((quads_crt_sva_8_376_296[80:54]),
          rec_quad_color_b_sva, or_tmp_328);
      rec_quad_color_g_sva_dfm <= MUX_v_27_2_2((quads_crt_sva_8_376_296[53:27]),
          rec_quad_color_g_sva, or_tmp_328);
      rec_quad_color_r_sva_dfm <= MUX_v_27_2_2((quads_crt_sva_8_376_296[26:0]), rec_quad_color_r_sva,
          or_tmp_328);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_hit_anything_sva_dfm <= 1'b0;
    end
    else if ( hit_wen & (fsm_output[2]) & for_stage_0_9 ) begin
      quad_hit_anything_sva_dfm <= quad_hit_anything_sva_dfm_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_normal_z_sva_dfm <= 26'b00000000000000000000000000;
      rec_quad_normal_y_sva_dfm <= 26'b00000000000000000000000000;
      rec_quad_normal_x_sva_dfm <= 26'b00000000000000000000000000;
    end
    else if ( rec_quad_normal_z_and_cse ) begin
      rec_quad_normal_z_sva_dfm <= MUX_v_26_2_2(quadInters_setfacenorm_run_qr_z_lpi_2_dfm_4_mx1w0,
          rec_quad_normal_z_sva, or_tmp_481);
      rec_quad_normal_y_sva_dfm <= MUX_v_26_2_2(quadInters_setfacenorm_run_qr_y_lpi_2_dfm_4_mx1w0,
          rec_quad_normal_y_sva, or_tmp_481);
      rec_quad_normal_x_sva_dfm <= MUX_v_26_2_2(quadInters_setfacenorm_run_qr_x_lpi_2_dfm_4_mx1w0,
          rec_quad_normal_x_sva, or_tmp_481);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_hit_loc_z_0_sva_dfm <= 1'b0;
      rec_quad_hit_loc_y_0_sva_dfm <= 1'b0;
      rec_quad_hit_loc_x_0_sva_dfm <= 1'b0;
    end
    else if ( rec_quad_hit_loc_z_and_cse ) begin
      rec_quad_hit_loc_z_0_sva_dfm <= MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_6_mx0w1,
          rec_quad_hit_loc_z_0_sva, or_tmp_490);
      rec_quad_hit_loc_y_0_sva_dfm <= MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_5_mx0w1,
          rec_quad_hit_loc_y_0_sva, or_tmp_490);
      rec_quad_hit_loc_x_0_sva_dfm <= MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_mx0w1,
          rec_quad_hit_loc_x_0_sva, or_tmp_490);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      add_run_ac_fixed_cctor_2_74_43_sva <= 32'b00000000000000000000000000000000;
      add_run_ac_fixed_cctor_1_74_43_sva <= 32'b00000000000000000000000000000000;
      add_run_ac_fixed_cctor_74_43_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( add_run_and_3_cse ) begin
      add_run_ac_fixed_cctor_2_74_43_sva <= add_run_ac_fixed_cctor_2_74_43_sva_mx1w0;
      add_run_ac_fixed_cctor_1_74_43_sva <= add_run_ac_fixed_cctor_1_74_43_sva_mx1w0;
      add_run_ac_fixed_cctor_74_43_sva <= add_run_ac_fixed_cctor_74_43_sva_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_run_lor_lpi_2_dfm <= 1'b0;
    end
    else if ( hit_wen & and_dcpl_54 & (fsm_output[3]) ) begin
      quadInters_run_lor_lpi_2_dfm <= quadInters_run_lor_lpi_2_dfm_mx0w1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_33_true_asn_1_itm_9 <= 1'b0;
    end
    else if ( hit_wen & (or_tmp_480 | or_tmp_481 | operator_33_true_asn_1_itm_9_mx0c2)
        ) begin
      operator_33_true_asn_1_itm_9 <= MUX1HOT_s_1_3_2(quadInters_run_quadInters_run_nor_4_cse_1,
          rec_quad_front_face_sva, operator_33_true_asn_1_itm_8, {or_tmp_480 , or_tmp_481
          , operator_33_true_asn_1_itm_9_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quads_crt_sva_8_110_108 <= 3'b000;
    end
    else if ( closest_so_far_and_cse & ((~ (fsm_output[5])) | rec_quad_mat_and_1_rgt)
        ) begin
      quads_crt_sva_8_110_108 <= MUX_v_3_2_2(rec_quad_mat_sva, (quads_crt_sva_7_110_0[110:108]),
          rec_quad_mat_and_1_rgt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_abs_21_21_1_xabs_xor_ftd_1 <= 20'b00000000000000000000;
      reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1 <= 20'b00000000000000000000;
      reg_ac_math_ac_abs_21_21_xabs_xor_ftd_1 <= 20'b00000000000000000000;
    end
    else if ( and_2744_cse ) begin
      reg_ac_math_ac_abs_21_21_1_xabs_xor_ftd_1 <= MUX_v_20_2_2((rec_quad_hit_loc_x_asn_ac_math_ac_abs_21_21_1_xabs_xor_itm_mx1w1_19_and_nl),
          (ac_math_ac_abs_21_21_1_xabs_xor_1_nl), ac_math_ac_abs_21_21_1_xabs_and_1_cse);
      reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1 <= MUX_v_20_2_2((rec_quad_hit_loc_y_asn_ac_math_ac_abs_21_21_2_xabs_xor_itm_mx1w1_19_and_nl),
          (ac_math_ac_abs_21_21_2_xabs_xor_1_nl), ac_math_ac_abs_21_21_1_xabs_and_1_cse);
      reg_ac_math_ac_abs_21_21_xabs_xor_ftd_1 <= MUX_v_20_2_2((rec_quad_hit_loc_z_asn_ac_math_ac_abs_21_21_xabs_xor_itm_mx1w1_19_and_nl),
          (ac_math_ac_abs_21_21_xabs_xor_1_nl), ac_math_ac_abs_21_21_1_xabs_and_1_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_run_lor_lpi_2_dfm_1 <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_8 <= 1'b0;
      quads_crt_sva_8_189_112 <= 78'b000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_8 <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_7 <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_5 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_6 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4
          <= 34'b0000000000000000000000000000000000;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_4 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_5 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3
          <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_4 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2
          <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_3 <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_1 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_st_2 <= 1'b0;
      quads_crt_sva_1_376_112 <= 265'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quadInters_run_land_lpi_2_dfm_st_1 <= 1'b0;
      quads_crt_sva_9_189_112 <= 78'b000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quadInters_run_lor_3_lpi_2_dfm_1 <= 1'b0;
      quadInters_run_land_lpi_2_dfm_9 <= 1'b0;
      quads_crt_sva_7_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      mult_run_asn_2_itm_1_74_30 <= 45'b000000000000000000000000000000000000000000000;
      quads_crt_sva_7_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quadInters_run_t_trunc_lpi_2_dfm_2_46 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_45 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_44 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_43 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_42 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_41 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_40 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_39 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_38 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_37 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_36 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_35 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_34 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_33 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_32 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_31 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_30 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_29 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_28 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_27 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_26 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_25 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_24 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_23 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_22 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_21 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_20 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_19 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_18 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_17 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_16 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_15 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_14 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_13 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_12 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_11 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_10 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_9 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_8 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_7 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_6 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_5 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_4 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_3 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_2 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_1 <= 1'b0;
      quadInters_run_t_trunc_lpi_2_dfm_2_0 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3
          <= 34'b0000000000000000000000000000000000;
      quads_crt_sva_7_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= 1'b0;
      operator_33_true_asn_1_itm_7 <= 1'b0;
      reg_quadInters_run_if_4_slc_quadInters_run_if_4_acc_27_svs_st_1_cse <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_9_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3
          <= 1'b0;
      quads_crt_sva_6_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_6_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2
          <= 34'b0000000000000000000000000000000000;
      quads_crt_sva_6_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_5_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_5_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_6 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_2
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0
          <= 22'b0000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1
          <= 34'b0000000000000000000000000000000000;
      quads_crt_sva_5_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_5 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_1
          <= 1'b0;
      quads_crt_sva_4_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_4_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_4_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_4 <= 1'b0;
      quads_crt_sva_3_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_3_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_3_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_3 <= 1'b0;
      quads_crt_sva_2_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_2_264_112 <= 153'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_1_110_0 <= 111'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      quads_crt_sva_2_376_296 <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_33_true_asn_1_itm_2 <= 1'b0;
      operator_33_true_asn_1_itm_1 <= 1'b0;
    end
    else if ( quadInters_run_oelse_and_1_cse ) begin
      quadInters_run_lor_lpi_2_dfm_1 <= quadInters_run_lor_lpi_2_dfm;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6;
      quadInters_run_land_lpi_2_dfm_8 <= quadInters_run_land_lpi_2_dfm_st_7;
      quads_crt_sva_8_189_112 <= quads_crt_sva_7_264_112[77:0];
      operator_33_true_asn_1_itm_8 <= operator_33_true_asn_1_itm_7;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_6 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_5;
      quadInters_run_land_lpi_2_dfm_st_7 <= quadInters_run_land_lpi_2_dfm_st_6;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_5 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_4;
      quadInters_run_land_lpi_2_dfm_st_6 <= quadInters_run_land_lpi_2_dfm_st_5;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_4 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3;
      quadInters_run_land_lpi_2_dfm_st_5 <= quadInters_run_land_lpi_2_dfm_st_4;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_3
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2;
      quadInters_run_land_lpi_2_dfm_st_4 <= quadInters_run_land_lpi_2_dfm_st_3;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_1;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_2 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_1;
      quadInters_run_land_lpi_2_dfm_st_3 <= quadInters_run_land_lpi_2_dfm_st_2;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_1 <= quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs;
      quadInters_run_land_lpi_2_dfm_st_2 <= quadInters_run_land_lpi_2_dfm_st_1;
      quads_crt_sva_1_376_112 <= quads_crt_sva[376:112];
      quadInters_run_land_lpi_2_dfm_st_1 <= quadInters_run_land_lpi_2_dfm;
      quads_crt_sva_9_189_112 <= quads_crt_sva_8_189_112;
      quadInters_run_lor_3_lpi_2_dfm_1 <= quadInters_run_lor_3_lpi_2_dfm;
      quadInters_run_land_lpi_2_dfm_9 <= quadInters_run_land_lpi_2_dfm_8;
      quads_crt_sva_7_110_0 <= quads_crt_sva_6_110_0;
      mult_run_asn_2_itm_1_74_30 <= mult_run_mul_cmp_z_oreg;
      quads_crt_sva_7_264_112 <= quads_crt_sva_6_264_112;
      quadInters_run_t_trunc_lpi_2_dfm_2_46 <= quadInters_run_t_trunc_lpi_2_dfm_1_46;
      quadInters_run_t_trunc_lpi_2_dfm_2_45 <= quadInters_run_t_trunc_lpi_2_dfm_1_45;
      quadInters_run_t_trunc_lpi_2_dfm_2_44 <= quadInters_run_t_trunc_lpi_2_dfm_1_44;
      quadInters_run_t_trunc_lpi_2_dfm_2_43 <= quadInters_run_t_trunc_lpi_2_dfm_1_43;
      quadInters_run_t_trunc_lpi_2_dfm_2_42 <= quadInters_run_t_trunc_lpi_2_dfm_1_42;
      quadInters_run_t_trunc_lpi_2_dfm_2_41 <= quadInters_run_t_trunc_lpi_2_dfm_1_41;
      quadInters_run_t_trunc_lpi_2_dfm_2_40 <= quadInters_run_t_trunc_lpi_2_dfm_1_40;
      quadInters_run_t_trunc_lpi_2_dfm_2_39 <= quadInters_run_t_trunc_lpi_2_dfm_1_39;
      quadInters_run_t_trunc_lpi_2_dfm_2_38 <= quadInters_run_t_trunc_lpi_2_dfm_1_38;
      quadInters_run_t_trunc_lpi_2_dfm_2_37 <= quadInters_run_t_trunc_lpi_2_dfm_1_37;
      quadInters_run_t_trunc_lpi_2_dfm_2_36 <= quadInters_run_t_trunc_lpi_2_dfm_1_36;
      quadInters_run_t_trunc_lpi_2_dfm_2_35 <= quadInters_run_t_trunc_lpi_2_dfm_1_35;
      quadInters_run_t_trunc_lpi_2_dfm_2_34 <= quadInters_run_t_trunc_lpi_2_dfm_1_34;
      quadInters_run_t_trunc_lpi_2_dfm_2_33 <= quadInters_run_t_trunc_lpi_2_dfm_1_33;
      quadInters_run_t_trunc_lpi_2_dfm_2_32 <= quadInters_run_t_trunc_lpi_2_dfm_1_32;
      quadInters_run_t_trunc_lpi_2_dfm_2_31 <= quadInters_run_t_trunc_lpi_2_dfm_1_31;
      quadInters_run_t_trunc_lpi_2_dfm_2_30 <= quadInters_run_t_trunc_lpi_2_dfm_1_30;
      quadInters_run_t_trunc_lpi_2_dfm_2_29 <= quadInters_run_t_trunc_lpi_2_dfm_1_29;
      quadInters_run_t_trunc_lpi_2_dfm_2_28 <= quadInters_run_t_trunc_lpi_2_dfm_1_28;
      quadInters_run_t_trunc_lpi_2_dfm_2_27 <= quadInters_run_t_trunc_lpi_2_dfm_1_27;
      quadInters_run_t_trunc_lpi_2_dfm_2_26 <= quadInters_run_t_trunc_lpi_2_dfm_1_26;
      quadInters_run_t_trunc_lpi_2_dfm_2_25 <= quadInters_run_t_trunc_lpi_2_dfm_1_25;
      quadInters_run_t_trunc_lpi_2_dfm_2_24 <= quadInters_run_t_trunc_lpi_2_dfm_1_24;
      quadInters_run_t_trunc_lpi_2_dfm_2_23 <= quadInters_run_t_trunc_lpi_2_dfm_1_23;
      quadInters_run_t_trunc_lpi_2_dfm_2_22 <= quadInters_run_t_trunc_lpi_2_dfm_1_22;
      quadInters_run_t_trunc_lpi_2_dfm_2_21 <= quadInters_run_t_trunc_lpi_2_dfm_1_21;
      quadInters_run_t_trunc_lpi_2_dfm_2_20 <= quadInters_run_t_trunc_lpi_2_dfm_1_20;
      quadInters_run_t_trunc_lpi_2_dfm_2_19 <= quadInters_run_t_trunc_lpi_2_dfm_1_19;
      quadInters_run_t_trunc_lpi_2_dfm_2_18 <= quadInters_run_t_trunc_lpi_2_dfm_1_18;
      quadInters_run_t_trunc_lpi_2_dfm_2_17 <= quadInters_run_t_trunc_lpi_2_dfm_1_17;
      quadInters_run_t_trunc_lpi_2_dfm_2_16 <= quadInters_run_t_trunc_lpi_2_dfm_1_16;
      quadInters_run_t_trunc_lpi_2_dfm_2_15 <= quadInters_run_t_trunc_lpi_2_dfm_1_15;
      quadInters_run_t_trunc_lpi_2_dfm_2_14 <= quadInters_run_t_trunc_lpi_2_dfm_1_14;
      quadInters_run_t_trunc_lpi_2_dfm_2_13 <= quadInters_run_t_trunc_lpi_2_dfm_1_13;
      quadInters_run_t_trunc_lpi_2_dfm_2_12 <= quadInters_run_t_trunc_lpi_2_dfm_1_12;
      quadInters_run_t_trunc_lpi_2_dfm_2_11 <= quadInters_run_t_trunc_lpi_2_dfm_1_11;
      quadInters_run_t_trunc_lpi_2_dfm_2_10 <= quadInters_run_t_trunc_lpi_2_dfm_1_10;
      quadInters_run_t_trunc_lpi_2_dfm_2_9 <= quadInters_run_t_trunc_lpi_2_dfm_1_9;
      quadInters_run_t_trunc_lpi_2_dfm_2_8 <= quadInters_run_t_trunc_lpi_2_dfm_1_8;
      quadInters_run_t_trunc_lpi_2_dfm_2_7 <= quadInters_run_t_trunc_lpi_2_dfm_1_7;
      quadInters_run_t_trunc_lpi_2_dfm_2_6 <= quadInters_run_t_trunc_lpi_2_dfm_1_6;
      quadInters_run_t_trunc_lpi_2_dfm_2_5 <= quadInters_run_t_trunc_lpi_2_dfm_1_5;
      quadInters_run_t_trunc_lpi_2_dfm_2_4 <= quadInters_run_t_trunc_lpi_2_dfm_1_4;
      quadInters_run_t_trunc_lpi_2_dfm_2_3 <= quadInters_run_t_trunc_lpi_2_dfm_1_3;
      quadInters_run_t_trunc_lpi_2_dfm_2_2 <= quadInters_run_t_trunc_lpi_2_dfm_1_2;
      quadInters_run_t_trunc_lpi_2_dfm_2_1 <= quadInters_run_t_trunc_lpi_2_dfm_1_1;
      quadInters_run_t_trunc_lpi_2_dfm_2_0 <= quadInters_run_t_trunc_lpi_2_dfm_1_0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ (z_out_6[33])), operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33])),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33])),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33])),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva[33])),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_2_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_3_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_4_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_1_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_5_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_33),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_33),
          operator_35_true_and_30_rgt);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_9_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_20_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33]),
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (z_out_6[33]), {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_18_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1[33]),
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33]),
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33]),
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_6_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_itm_1,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_33_itm,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_3_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_33_itm,
          {operator_35_true_and_30_rgt , operator_35_true_and_31_rgt , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33
          <= z_out_4[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2;
      quads_crt_sva_7_376_296 <= quads_crt_sva_6_376_296;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      operator_33_true_asn_1_itm_7 <= operator_33_true_asn_1_itm_6;
      reg_quadInters_run_if_4_slc_quadInters_run_if_4_acc_27_svs_st_1_cse <= readslicef_28_1_27((quadInters_run_if_4_acc_nl));
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_33_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[33];
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_33_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= z_out_7[33];
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_9_psp_33_itm_1
          <= reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_33_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_33_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_itm_1
          <= operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_3
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_2;
      quads_crt_sva_6_110_0 <= quads_crt_sva_5_110_0;
      quads_crt_sva_6_264_112 <= quads_crt_sva_5_264_112;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1;
      quads_crt_sva_6_376_296 <= quads_crt_sva_5_376_296;
      quads_crt_sva_5_110_0 <= quads_crt_sva_4_110_0;
      quads_crt_sva_5_264_112 <= quads_crt_sva_4_264_112;
      operator_33_true_asn_1_itm_6 <= operator_33_true_asn_1_itm_5;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_26_sva_1[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= z_out_9[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= z_out_10[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_2
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0
          <= quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24[21:0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm;
      quads_crt_sva_5_376_296 <= quads_crt_sva_4_376_296;
      operator_33_true_asn_1_itm_5 <= operator_33_true_asn_1_itm_4;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_1
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs;
      quads_crt_sva_4_110_0 <= quads_crt_sva_3_110_0;
      quads_crt_sva_4_264_112 <= quads_crt_sva_3_264_112;
      quads_crt_sva_4_376_296 <= quads_crt_sva_3_376_296;
      operator_33_true_asn_1_itm_4 <= operator_33_true_asn_1_itm_3;
      quads_crt_sva_3_110_0 <= quads_crt_sva_2_110_0;
      quads_crt_sva_3_264_112 <= quads_crt_sva_2_264_112;
      quads_crt_sva_3_376_296 <= quads_crt_sva_2_376_296;
      operator_33_true_asn_1_itm_3 <= operator_33_true_asn_1_itm_2;
      quads_crt_sva_2_110_0 <= quads_crt_sva_1_110_0;
      quads_crt_sva_2_264_112 <= quads_crt_sva_1_376_112[152:0];
      quads_crt_sva_1_110_0 <= quads_crt_sva[110:0];
      quads_crt_sva_2_376_296 <= quads_crt_sva_1_376_112[264:184];
      operator_33_true_asn_1_itm_2 <= operator_33_true_asn_1_itm_1;
      operator_33_true_asn_1_itm_1 <= operator_33_true_asn_1_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_hit_loc_z_20_1_sva <= 20'b00000000000000000000;
      rec_quad_hit_loc_y_20_1_sva <= 20'b00000000000000000000;
      rec_quad_hit_loc_x_20_1_sva <= 20'b00000000000000000000;
    end
    else if ( and_2754_cse ) begin
      rec_quad_hit_loc_z_20_1_sva <= MUX_v_20_2_2(20'b00000000000000000000, quadInters_run_quadInters_run_and_6_mx0w2,
          (not_676_nl));
      rec_quad_hit_loc_y_20_1_sva <= MUX_v_20_2_2(20'b00000000000000000000, quadInters_run_quadInters_run_and_4_mx0w2,
          (not_674_nl));
      rec_quad_hit_loc_x_20_1_sva <= MUX_v_20_2_2(20'b00000000000000000000, quadInters_run_quadInters_run_and_2_mx0w2,
          (not_672_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_color_b_sva <= 27'b000000000000000000000000000;
      rec_quad_color_g_sva <= 27'b000000000000000000000000000;
      rec_quad_color_r_sva <= 27'b000000000000000000000000000;
      rec_quad_mat_sva <= 3'b000;
    end
    else if ( and_2778_cse ) begin
      rec_quad_color_b_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, (quads_crt_sva_8_376_296[80:54]),
          (rec_quad_color_b_not_nl));
      rec_quad_color_g_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, (quads_crt_sva_8_376_296[53:27]),
          (rec_quad_color_g_not_nl));
      rec_quad_color_r_sva <= MUX_v_27_2_2(27'b000000000000000000000000000, (quads_crt_sva_8_376_296[26:0]),
          (rec_quad_color_r_not_nl));
      rec_quad_mat_sva <= MUX_v_3_2_2(3'b000, quads_crt_sva_8_110_108, (rec_quad_mat_not_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56 <= 2'b00;
    end
    else if ( ((quadInters_run_if_1_acc_itm_34 & (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs)
        & (fsm_output[3])) | (fsm_output[5:4]!=2'b00)) & hit_wen ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_1_57_56 <= quadInters_denom_dot_run_mux1h_5_rgt[33:32];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24 <= 32'b00000000000000000000000000000000;
    end
    else if ( ((~((~((quadInters_run_if_1_acc_itm_34 & (fsm_output[3])) | (fsm_output[4])))
        | quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs)) | (fsm_output[5]))
        & hit_wen ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_1_55_24 <= quadInters_denom_dot_run_mux1h_5_rgt[31:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_i_5_0_sva_4_0 <= 5'b00000;
    end
    else if ( (((fsm_output[5:3]==3'b000) & for_stage_0_1) | (fsm_output[6]) | (fsm_output[0])
        | (fsm_output[1])) & hit_wen ) begin
      for_i_5_0_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_1[4:0]), (not_671_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quad_max_sva <= 11'b00000000000;
    end
    else if ( hit_wen & (~ or_tmp_691) ) begin
      quad_max_sva <= quad_max_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rec_quad_normal_z_sva <= 26'b00000000000000000000000000;
      rec_quad_normal_y_sva <= 26'b00000000000000000000000000;
      rec_quad_normal_x_sva <= 26'b00000000000000000000000000;
    end
    else if ( and_2828_cse ) begin
      rec_quad_normal_z_sva <= MUX_v_26_2_2(26'b00000000000000000000000000, quadInters_setfacenorm_run_qr_z_lpi_2_dfm_4_mx1w0,
          (rec_quad_normal_z_not_nl));
      rec_quad_normal_y_sva <= MUX_v_26_2_2(26'b00000000000000000000000000, quadInters_setfacenorm_run_qr_y_lpi_2_dfm_4_mx1w0,
          (rec_quad_normal_y_not_nl));
      rec_quad_normal_x_sva <= MUX_v_26_2_2(26'b00000000000000000000000000, quadInters_setfacenorm_run_qr_x_lpi_2_dfm_4_mx1w0,
          (rec_quad_normal_x_not_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_setfacenorm_run_qr_z_lpi_2 <= 26'b00000000000000000000000000;
      quadInters_setfacenorm_run_qr_y_lpi_2 <= 26'b00000000000000000000000000;
      quadInters_setfacenorm_run_qr_x_lpi_2 <= 26'b00000000000000000000000000;
    end
    else if ( and_2843_cse ) begin
      quadInters_setfacenorm_run_qr_z_lpi_2 <= quadInters_setfacenorm_run_qr_z_lpi_2_dfm_4_mx1w0;
      quadInters_setfacenorm_run_qr_y_lpi_2 <= quadInters_setfacenorm_run_qr_y_lpi_2_dfm_4_mx1w0;
      quadInters_setfacenorm_run_qr_x_lpi_2 <= quadInters_setfacenorm_run_qr_x_lpi_2_dfm_4_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_run_lor_lpi_2_dfm_2 <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_1_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_33_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_33_itm
          <= 1'b0;
    end
    else if ( quadInters_run_oelse_and_2_cse ) begin
      quadInters_run_lor_lpi_2_dfm_2 <= MUX_s_1_2_2(quadInters_run_lor_lpi_2_dfm_mx0w1,
          quadInters_run_lor_lpi_2_dfm_1, fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_1_itm_1
          <= MUX_s_1_2_2((z_out_7[33]), (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[1]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]),
          (add_run_ac_fixed_cctor_1_74_43_sva[31]), fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((z_out_12[34]), (add_run_ac_fixed_cctor_2_74_43_sva[31]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((z_out_11[34]), (add_run_ac_fixed_cctor_74_43_sva[31]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_psp_sva_1[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[0]),
          fsm_output[5]);
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_1_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1[33]),
          reg_quadInters_run_if_4_slc_quadInters_run_if_4_acc_27_svs_st_1_cse, fsm_output[5]);
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_33_itm
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33,
          quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7, fsm_output[5]);
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_33_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[33]),
          quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_7, fsm_output[5]);
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_33_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[33]),
          reg_quadInters_run_if_4_slc_quadInters_run_if_4_acc_27_svs_st_1_cse, fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
    end
    else if ( operator_35_true_and_59_cse ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_4_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {(fsm_output[4]) , operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_4_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_6_psp_sva_1[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {(fsm_output[4]) , operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_4_2((z_out_5[33]), (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {(fsm_output[4]) , operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_4_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_5_psp_sva_1[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {(fsm_output[4]) , operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1
          <= MUX1HOT_s_1_4_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm_1,
          {(fsm_output[4]) , operator_35_true_and_30_rgt , operator_35_true_and_31_rgt
          , operator_35_true_and_32_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((z_out_13[34]), div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2,
          fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_stage_0_1 <= 1'b0;
      for_stage_0_2 <= 1'b0;
      for_stage_0_3 <= 1'b0;
      for_stage_0_4 <= 1'b0;
      for_stage_0_5 <= 1'b0;
      for_stage_0_6 <= 1'b0;
      for_stage_0_7 <= 1'b0;
      for_stage_0_8 <= 1'b0;
      for_stage_0_9 <= 1'b0;
    end
    else if ( for_and_1_cse ) begin
      for_stage_0_1 <= for_stage_0 | (fsm_output[1]);
      for_stage_0_2 <= for_stage_0_1 & (~ (fsm_output[1]));
      for_stage_0_3 <= for_stage_0_2 & (~ (fsm_output[1]));
      for_stage_0_4 <= for_stage_0_3 & (~ (fsm_output[1]));
      for_stage_0_5 <= for_stage_0_4 & (~ (fsm_output[1]));
      for_stage_0_6 <= for_stage_0_5 & (~ (fsm_output[1]));
      for_stage_0_7 <= for_stage_0_6 & (~ (fsm_output[1]));
      for_stage_0_8 <= for_stage_0_7 & (~ (fsm_output[1]));
      for_stage_0_9 <= for_stage_0_8 & (~ (fsm_output[1]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_47_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_46_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
    end
    else if ( operator_35_true_and_100_cse ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_67_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ (z_out_6[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_66_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_65_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_32_psp_sva_1[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_31_psp_sva_1[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_56_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_55_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_54_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_53_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_20_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_52_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_51_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_18_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_50_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_49_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_48_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_47_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_46_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= ~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= 1'b0;
    end
    else if ( operator_35_true_and_135_cse ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_33_1_itm,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[33]),
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_11_psp_sva_1[33]),
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_12_psp_sva_1[33]),
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          (z_out_7[33]), operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          operator_35_true_and_282_cse);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm
          <= MUX_s_1_2_2((~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_2),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm,
          operator_35_true_and_282_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_2_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_3_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_4_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_6_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      quadInters_run_lor_3_lpi_2_dfm <= 1'b0;
      for_hitWorld_lpi_2_dfm_2 <= 1'b0;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs <= 1'b0;
      quadInters_run_land_lpi_2_dfm <= 1'b0;
      quads_crt_sva <= 377'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_18_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= 1'b0;
      operator_33_true_asn_1_itm <= 1'b0;
    end
    else if ( div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_cse
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_2_itm_1
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33,
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[2]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_3_itm_1
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[3]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_4_itm_1
          <= MUX_s_1_2_2((z_out_5[33]), (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[4]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_6_itm_1
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[6]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_46_lpi_2_dfm_mx0[0]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= MUX_s_1_2_2((z_out_10[34]), (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_68_lpi_2_dfm_mx0[0]),
          fsm_output[5]);
      quadInters_run_lor_3_lpi_2_dfm <= quadInters_run_if_5_quadInters_run_if_5_or_2_tmp;
      for_hitWorld_lpi_2_dfm_2 <= for_hitWorld_lpi_2_dfm_3;
      quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs <= readslicef_35_1_34((quadInters_run_if_2_acc_nl));
      quadInters_run_land_lpi_2_dfm <= (quads_rsci_idat_mxwt[111]) & (ray_temp_in_crt_sva[165]);
      quads_crt_sva <= quads_rsci_idat_mxwt;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_33_itm
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_18_psp_sva_33
          <= z_out_5[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_16_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_15_psp_sva_1[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_31_sva_1[34];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_30_sva_1[34];
      operator_33_true_asn_1_itm <= or_343_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_5_itm_1
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_20_psp_sva_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33
          <= 1'b0;
    end
    else if ( div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_and_3_cse
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_5_itm_1
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[5]),
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_23_psp_sva_mx0w0[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_22_psp_sva_mx0w0[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_21_psp_sva_mx0w0[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_20_psp_sva_33
          <= z_out_7[33];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1[33];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_itm
          <= 34'b0000000000000000000000000000000000;
    end
    else if ( hit_wen & (((~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs)
        & (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0[34])
        & (fsm_output[5])) | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_6_rgt)
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_itm
          <= MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_6_rgt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33
          <= 1'b0;
    end
    else if ( or_1462_cse & hit_wen ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_11_rgt[33];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_32_0
          <= 33'b000000000000000000000000000000000;
    end
    else if ( ((fsm_output[5:2]!=4'b0000)) & hit_wen ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_32_0
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_11_rgt[32:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st
          <= 1'b0;
    end
    else if ( div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_5_cse
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva
          <= MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
          fsm_output[5]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_st
          <= MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_mx1w0,
          for_hitWorld_lpi_2_dfm_2, fsm_output[5]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_abs_58_58_xabs_xor_itm <= 58'b0000000000000000000000000000000000000000000000000000000000;
    end
    else if ( hit_wen & (~((fsm_output[3]) | (quadInters_run_land_lpi_2_dfm & (fsm_output[4]))
        | quadInters_denom_dot_run_and_5_rgt)) ) begin
      ac_math_ac_abs_58_58_xabs_xor_itm <= MUX_v_58_2_2((quadInters_denom_dot_run_acc_2_nl),
          (ac_math_ac_abs_58_58_xabs_xor_nl), quadInters_denom_dot_run_and_4_rgt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_33_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_33_itm
          <= 1'b0;
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_33_itm
          <= 1'b0;
    end
    else if ( operator_35_true_and_185_cse ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= MUX1HOT_s_1_3_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_33,
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_33_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm
          <= MUX1HOT_s_1_3_2((z_out_6[33]), (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm_1),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_34_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_33_itm
          <= MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_sva_mx0w1[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_45_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_33_itm
          <= MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_46_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_33_itm
          <= MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1[33]),
          (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_14_psp_sva_1_33),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_47_operator_80_false_operator_80_false_operator_35_true_not_1_itm,
          {(fsm_output[4]) , operator_35_true_and_16_rgt , operator_35_true_and_31_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva
          <= 35'b00000000000000000000000000000000000;
    end
    else if ( hit_wen & (~((fsm_output[3]) | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_1_cse
        | (quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs & (fsm_output[5]))))
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva
          <= MUX1HOT_v_35_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_8_sva_mx2w0,
          {(fsm_output[2]) , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_rgt
          , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl)});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      setfacenorm_dot_run_acc_2_itm <= 60'b000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( hit_wen & (~(or_dcpl_79 | (quadInters_run_lor_3_lpi_2_dfm & (fsm_output[5]))))
        ) begin
      setfacenorm_dot_run_acc_2_itm <= MUX_v_60_2_2(z_out, quadInters_denom_dot_run_mul_1_cmp_z_oreg,
          setfacenorm_dot_run_and_1_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg <= 21'b000000000000000000000;
      reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg <= 21'b000000000000000000000;
      reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg <= 21'b000000000000000000000;
    end
    else if ( and_2862_cse ) begin
      reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg <= quadInters_sub_run_mux_rgt[20:0];
      reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg <= quadInters_sub_run_mux_1_rgt[20:0];
      reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg <= quadInters_sub_run_mux_2_rgt[20:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mult_run_asn_1_itm_42_30 <= 13'b0000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd
          <= 1'b0;
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd
          <= 1'b0;
    end
    else if ( and_2865_cse ) begin
      mult_run_asn_1_itm_42_30 <= mult_run_mul_cmp_z_oreg[12:0];
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_42_psp_sva_33
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_65_rgt[33];
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_sva_1[33]),
          (z_out_2[33]), fsm_output[4]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_ftd
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_37_psp_sva_1[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_26_psp_sva_mx0w2[33]),
          fsm_output[4]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_ftd
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_38_psp_sva_1[33]),
          (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[33]),
          fsm_output[4]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_28_psp_ftd
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_39_psp_sva_1[33]),
          (z_out_6[33]), fsm_output[4]);
      reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_30_psp_ftd
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_40_psp_sva_1[33]),
          (z_out_3[33]), fsm_output[4]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33
          <= 1'b0;
    end
    else if ( (fsm_output[4:3]==2'b00) & hit_wen ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33
          <= z_out_2[33];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_57_24 <= 34'b0000000000000000000000000000000000;
    end
    else if ( (fsm_output[4]) & (~ quadInters_run_land_lpi_2_dfm) & hit_wen ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_57_24 <= quadInters_denom_dot_run_mul_2_cmp_1_z_oreg[57:24];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_23_0 <= 24'b000000000000000000000000;
    end
    else if ( (~((fsm_output[4]) & quadInters_run_land_lpi_2_dfm)) & hit_wen ) begin
      quadInters_denom_dot_run_ac_fixed_cctor_sva_23_0 <= quadInters_denom_dot_run_mul_2_cmp_1_z_oreg[23:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm
          <= 34'b0000000000000000000000000000000000;
    end
    else if ( hit_wen & (((~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs)
        & quadInters_run_mux_593_tmp_33 & (~ (fsm_output[4]))) | div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_and_rgt)
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm
          <= MUX_v_34_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl),
          ({1'b0 , quadInters_run_rounded_denom_lpi_2_dfm_mx0_32_0}), div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qelse_and_rgt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm
          <= 34'b0000000000000000000000000000000000;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_45
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_44
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_43
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_3
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_42
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_4
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_41
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_5
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_40
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_6
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_39
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_7
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_38
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_8
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_37
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_9
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_36
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_35
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_34
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_33
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_32
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_31
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_30
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_29
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_28
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_27
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_26
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_25
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_21
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_24
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_22
          <= 1'b0;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_23
          <= 1'b0;
    end
    else if ( div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_cse
        ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva
          <= div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1;
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_lpi_2_dfm
          <= MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_4,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1[33]);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[46]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_21_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_45
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[45]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_22_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_44
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[44]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_23_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_43
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[43]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_24_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_3
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[3]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_64_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_42
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[42]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_25_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_4
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[4]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_63_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_41
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[41]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_26_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_5
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[5]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_62_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_40
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[40]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_27_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_6
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[6]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_39
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[39]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_28_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_7
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[7]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_60_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_38
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[38]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_29_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_8
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[8]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_37
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[37]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_30_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_9
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[9]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_58_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_36
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[36]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_31_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_35
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[35]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_57_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_34
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[34]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_59_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_33
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[33]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_61_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_32
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[32]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_31
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[31]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_36_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_30
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[30]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_37_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_29
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[29]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_38_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_28
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[28]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_39_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_27
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[27]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_40_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_26
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[26]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_41_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_25
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[25]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_42_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_21
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[21]),
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_33_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_24
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[24]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_43_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_22
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[22]),
          operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_25_psp_33_itm,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_23
          <= MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[23]),
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_44_operator_80_false_operator_80_false_operator_35_true_not_1_itm_1,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_57_lpi_2_dfm
          <= 34'b0000000000000000000000000000000000;
    end
    else if ( hit_wen & for_stage_0_5 & (~ quadInters_run_land_lpi_2_dfm_st_4) &
        (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs_st_3) ) begin
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_57_lpi_2_dfm
          <= MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_3,
          div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_24_psp_sva_1[33]);
    end
  end
  assign quadInters_cross_u_run_mul_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[59:48]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg
      , (add_run_ac_fixed_cctor_2_74_43_sva[8:0]) , (mult_run_asn_2_itm_1_74_30[12:0])})));
  assign quadInters_cross_u_run_mul_1_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[71:60]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg
      , (add_run_ac_fixed_cctor_1_74_43_sva[8:0]) , mult_run_asn_1_itm_42_30})));
  assign nl_quadInters_cross_u_run_acc_nl = (quadInters_cross_u_run_mul_nl) - (quadInters_cross_u_run_mul_1_nl);
  assign quadInters_cross_u_run_acc_nl = nl_quadInters_cross_u_run_acc_nl[56:0];
  assign quadInters_cross_u_run_mul_4_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[47:36]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg
      , (add_run_ac_fixed_cctor_1_74_43_sva[8:0]) , mult_run_asn_1_itm_42_30})));
  assign quadInters_cross_u_run_mul_5_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[59:48]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg
      , (add_run_ac_fixed_cctor_74_43_sva[8:0]) , quadInters_at_run_mult_result_x_74_30_sva_12_0})));
  assign nl_quadInters_cross_u_run_acc_2_nl = (quadInters_cross_u_run_mul_4_nl) -
      (quadInters_cross_u_run_mul_5_nl);
  assign quadInters_cross_u_run_acc_2_nl = nl_quadInters_cross_u_run_acc_2_nl[56:0];
  assign quadInters_cross_v_run_mul_4_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg , (add_run_ac_fixed_cctor_74_43_sva[8:0])
      , quadInters_at_run_mult_result_x_74_30_sva_12_0})) * $signed((quads_crt_sva_7_110_0[95:84])));
  assign quadInters_cross_v_run_mul_5_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg , (add_run_ac_fixed_cctor_1_74_43_sva[8:0])
      , mult_run_asn_1_itm_42_30})) * $signed((quads_crt_sva_7_110_0[83:72])));
  assign nl_quadInters_cross_v_run_acc_2_nl = (quadInters_cross_v_run_mul_4_nl) -
      (quadInters_cross_v_run_mul_5_nl);
  assign quadInters_cross_v_run_acc_2_nl = nl_quadInters_cross_v_run_acc_2_nl[56:0];
  assign quadInters_cross_v_run_mul_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg , (add_run_ac_fixed_cctor_1_74_43_sva[8:0])
      , mult_run_asn_1_itm_42_30})) * $signed((quads_crt_sva_7_110_0[107:96])));
  assign quadInters_cross_v_run_mul_1_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg , (add_run_ac_fixed_cctor_2_74_43_sva[8:0])
      , (mult_run_asn_2_itm_1_74_30[12:0])})) * $signed((quads_crt_sva_7_110_0[95:84])));
  assign nl_quadInters_cross_v_run_acc_nl = (quadInters_cross_v_run_mul_nl) - (quadInters_cross_v_run_mul_1_nl);
  assign quadInters_cross_v_run_acc_nl = nl_quadInters_cross_v_run_acc_nl[56:0];
  assign quadInters_cross_u_run_mul_2_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[71:60]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg
      , (add_run_ac_fixed_cctor_74_43_sva[8:0]) , quadInters_at_run_mult_result_x_74_30_sva_12_0})));
  assign quadInters_cross_u_run_mul_3_nl = conv_s2u_57_57($signed((quads_crt_sva_7_110_0[47:36]))
      * $signed(({reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg , reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg
      , (add_run_ac_fixed_cctor_2_74_43_sva[8:0]) , (mult_run_asn_2_itm_1_74_30[12:0])})));
  assign nl_quadInters_cross_u_run_acc_1_nl = (quadInters_cross_u_run_mul_2_nl) -
      (quadInters_cross_u_run_mul_3_nl);
  assign quadInters_cross_u_run_acc_1_nl = nl_quadInters_cross_u_run_acc_1_nl[56:0];
  assign quad_hit_anything_mux_48_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_46, closest_so_far_sva_46,
      or_tmp_531);
  assign quad_hit_anything_mux_47_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_0, closest_so_far_sva_0,
      or_tmp_531);
  assign quad_hit_anything_mux_46_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_45, closest_so_far_sva_45,
      or_tmp_531);
  assign quad_hit_anything_mux_45_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_1, closest_so_far_sva_1,
      or_tmp_531);
  assign quad_hit_anything_mux_44_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_44, closest_so_far_sva_44,
      or_tmp_531);
  assign quad_hit_anything_mux_43_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_2, closest_so_far_sva_2,
      or_tmp_531);
  assign quad_hit_anything_mux_42_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_43, closest_so_far_sva_43,
      or_tmp_531);
  assign quad_hit_anything_mux_41_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_3, closest_so_far_sva_3,
      or_tmp_531);
  assign quad_hit_anything_mux_40_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_42, closest_so_far_sva_42,
      or_tmp_531);
  assign quad_hit_anything_mux_39_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_4, closest_so_far_sva_4,
      or_tmp_531);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_4_nl
      = MUX_s_1_2_2(closest_so_far_sva_dfm_3_41, closest_so_far_sva_41, or_tmp_531);
  assign quad_hit_anything_mux_38_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_5, closest_so_far_sva_5,
      or_tmp_531);
  assign quad_hit_anything_mux_37_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_40, closest_so_far_sva_40,
      or_tmp_531);
  assign quad_hit_anything_mux_36_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_6, closest_so_far_sva_6,
      or_tmp_531);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_3_nl
      = MUX_s_1_2_2(closest_so_far_sva_dfm_3_39, closest_so_far_sva_39, or_tmp_531);
  assign quad_hit_anything_mux_35_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_7, closest_so_far_sva_7,
      or_tmp_531);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_2_nl
      = MUX_s_1_2_2(closest_so_far_sva_dfm_3_38, closest_so_far_sva_38, or_tmp_531);
  assign quad_hit_anything_mux_34_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_8, closest_so_far_sva_8,
      or_tmp_531);
  assign quad_hit_anything_mux_33_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_37, closest_so_far_sva_37,
      or_tmp_531);
  assign quad_hit_anything_mux_32_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_9, closest_so_far_sva_9,
      or_tmp_531);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_1_nl
      = MUX_s_1_2_2(closest_so_far_sva_dfm_3_36, closest_so_far_sva_36, or_tmp_531);
  assign quad_hit_anything_mux_31_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_10, closest_so_far_sva_10,
      or_tmp_531);
  assign quad_hit_anything_mux_30_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_35, closest_so_far_sva_35,
      or_tmp_531);
  assign quad_hit_anything_mux_29_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_11, closest_so_far_sva_11,
      or_tmp_531);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_rem_oelse_mux_nl
      = MUX_s_1_2_2(closest_so_far_sva_dfm_3_34, closest_so_far_sva_34, or_tmp_531);
  assign quad_hit_anything_mux_28_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_12, closest_so_far_sva_12,
      or_tmp_531);
  assign quad_hit_anything_mux_27_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_33, closest_so_far_sva_33,
      or_tmp_531);
  assign quad_hit_anything_mux_26_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_13, closest_so_far_sva_13,
      or_tmp_531);
  assign quad_hit_anything_mux_25_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_32, closest_so_far_sva_32,
      or_tmp_531);
  assign quad_hit_anything_mux_24_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_14, closest_so_far_sva_14,
      or_tmp_531);
  assign quad_hit_anything_mux_23_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_31, closest_so_far_sva_31,
      or_tmp_531);
  assign quad_hit_anything_mux_22_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_15, closest_so_far_sva_15,
      or_tmp_531);
  assign quad_hit_anything_mux_21_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_30, closest_so_far_sva_30,
      or_tmp_531);
  assign quad_hit_anything_mux_20_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_16, closest_so_far_sva_16,
      or_tmp_531);
  assign quad_hit_anything_mux_19_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_29, closest_so_far_sva_29,
      or_tmp_531);
  assign quad_hit_anything_mux_18_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_17, closest_so_far_sva_17,
      or_tmp_531);
  assign quad_hit_anything_mux_17_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_28, closest_so_far_sva_28,
      or_tmp_531);
  assign quad_hit_anything_mux_16_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_18, closest_so_far_sva_18,
      or_tmp_531);
  assign quad_hit_anything_mux_15_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_27, closest_so_far_sva_27,
      or_tmp_531);
  assign quad_hit_anything_mux_14_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_19, closest_so_far_sva_19,
      or_tmp_531);
  assign quad_hit_anything_mux_13_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_26, closest_so_far_sva_26,
      or_tmp_531);
  assign quad_hit_anything_mux_12_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_20, closest_so_far_sva_20,
      or_tmp_531);
  assign quad_hit_anything_mux_11_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_25, closest_so_far_sva_25,
      or_tmp_531);
  assign quad_hit_anything_mux_10_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_21, closest_so_far_sva_21,
      or_tmp_531);
  assign quad_hit_anything_mux_9_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_24, closest_so_far_sva_24,
      or_tmp_531);
  assign quad_hit_anything_mux_8_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_22, closest_so_far_sva_22,
      or_tmp_531);
  assign quad_hit_anything_mux_7_nl = MUX_s_1_2_2(closest_so_far_sva_dfm_3_23, closest_so_far_sva_23,
      or_tmp_531);
  assign quad_hit_anything_mux_6_nl = MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_6_mx0w1,
      rec_quad_hit_loc_z_0_sva, or_tmp_673);
  assign quad_hit_anything_mux_5_nl = MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_5_mx0w1,
      rec_quad_hit_loc_y_0_sva, or_tmp_673);
  assign quad_hit_anything_mux_4_nl = MUX_s_1_2_2(quadInters_run_quadInters_run_quadInters_run_nor_mx0w1,
      rec_quad_hit_loc_x_0_sva, or_tmp_673);
  assign quad_hit_anything_mux_2_nl = MUX_s_1_2_2(quad_hit_anything_sva_dfm_mx0w0,
      quad_hit_anything_sva, or_dcpl_95);
  assign quad_hit_anything_mux_nl = MUX_s_1_2_2((quad_hit_anything_mux_2_nl), quad_hit_anything_sva,
      and_1128_cse);
  assign quad_hit_anything_mux_3_nl = MUX_s_1_2_2(rec_quad_front_face_sva, quadInters_run_quadInters_run_nor_4_cse_1,
      and_1706_cse);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_5_nl
      = (z_out_8[34]) & div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_m1c;
  assign quad_hit_anything_mux1h_58_nl = MUX1HOT_s_1_3_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_mx1w0,
      for_stage_0_9, {div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_or_rgt
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_and_rgt
      , (fsm_output[5])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_78_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_46_psp_sva_1[33]));
  assign operator_35_true_mux_172_nl = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_else_acc_itm_59_13[20]),
      operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_33_itm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_if_xnor_svs_4);
  assign mux_125_nl = MUX_v_20_2_2(quadInters_run_quadInters_run_and_2_mx0w2, rec_quad_hit_loc_x_20_1_sva,
      or_tmp_490);
  assign not_nl = ~ (fsm_output[0]);
  assign rec_quad_hit_loc_x_asn_ac_math_ac_abs_21_21_1_xabs_xor_itm_mx1w1_19_and_nl
      = MUX_v_20_2_2(20'b00000000000000000000, (mux_125_nl), (not_nl));
  assign ac_math_ac_abs_21_21_1_xabs_xor_1_nl = (signext_20_1(reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg[20]))
      ^ (reg_quadInters_sub_run_ac_fixed_cctor_1_44_22_1_reg[19:0]);
  assign mux_124_nl = MUX_v_20_2_2(quadInters_run_quadInters_run_and_4_mx0w2, rec_quad_hit_loc_y_20_1_sva,
      or_tmp_490);
  assign not_669_nl = ~ (fsm_output[0]);
  assign rec_quad_hit_loc_y_asn_ac_math_ac_abs_21_21_2_xabs_xor_itm_mx1w1_19_and_nl
      = MUX_v_20_2_2(20'b00000000000000000000, (mux_124_nl), (not_669_nl));
  assign ac_math_ac_abs_21_21_2_xabs_xor_1_nl = (signext_20_1(reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg[20]))
      ^ (reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg[19:0]);
  assign mux_123_nl = MUX_v_20_2_2(quadInters_run_quadInters_run_and_6_mx0w2, rec_quad_hit_loc_z_20_1_sva,
      or_tmp_490);
  assign not_670_nl = ~ (fsm_output[0]);
  assign rec_quad_hit_loc_z_asn_ac_math_ac_abs_21_21_xabs_xor_itm_mx1w1_19_and_nl
      = MUX_v_20_2_2(20'b00000000000000000000, (mux_123_nl), (not_670_nl));
  assign ac_math_ac_abs_21_21_xabs_xor_1_nl = (signext_20_1(reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg[20]))
      ^ (reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg[19:0]);
  assign nl_quadInters_run_if_4_acc_nl = conv_s2u_27_28({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_else_Q_60_14_lpi_2_dfm_46
      , quadInters_run_t_trunc_lpi_2_dfm_45_1 , quadInters_run_t_trunc_lpi_2_dfm_44_1
      , quadInters_run_t_trunc_lpi_2_dfm_43_1 , quadInters_run_t_trunc_lpi_2_dfm_42_1
      , quadInters_run_t_trunc_lpi_2_dfm_41_1 , quadInters_run_t_trunc_lpi_2_dfm_40_1
      , quadInters_run_t_trunc_lpi_2_dfm_39_1 , quadInters_run_t_trunc_lpi_2_dfm_38_1
      , quadInters_run_t_trunc_lpi_2_dfm_37_1 , quadInters_run_t_trunc_lpi_2_dfm_36_1
      , quadInters_run_t_trunc_lpi_2_dfm_35_1 , quadInters_run_t_trunc_lpi_2_dfm_34_1
      , quadInters_run_t_trunc_lpi_2_dfm_33_1 , quadInters_run_t_trunc_lpi_2_dfm_32_1
      , quadInters_run_t_trunc_lpi_2_dfm_31_1 , quadInters_run_t_trunc_lpi_2_dfm_30_1
      , quadInters_run_t_trunc_lpi_2_dfm_29_1 , quadInters_run_t_trunc_lpi_2_dfm_28_1
      , quadInters_run_t_trunc_lpi_2_dfm_27_1 , quadInters_run_t_trunc_lpi_2_dfm_26_1
      , quadInters_run_t_trunc_lpi_2_dfm_25_1 , quadInters_run_t_trunc_lpi_2_dfm_24_1
      , quadInters_run_t_trunc_lpi_2_dfm_23_1 , quadInters_run_t_trunc_lpi_2_dfm_22_1
      , quadInters_run_t_trunc_lpi_2_dfm_21_1 , quadInters_run_t_trunc_lpi_2_dfm_20_1})
      + 28'b1111111111111111111111111111;
  assign quadInters_run_if_4_acc_nl = nl_quadInters_run_if_4_acc_nl[27:0];
  assign not_676_nl = ~ or_tmp_529;
  assign not_674_nl = ~ or_tmp_529;
  assign not_672_nl = ~ or_tmp_529;
  assign rec_quad_color_b_not_nl = ~ or_tmp_529;
  assign rec_quad_color_g_not_nl = ~ or_tmp_529;
  assign rec_quad_color_r_not_nl = ~ or_tmp_529;
  assign rec_quad_mat_not_nl = ~ or_tmp_529;
  assign not_671_nl = ~ or_tmp_529;
  assign rec_quad_normal_z_not_nl = ~ or_tmp_529;
  assign rec_quad_normal_y_not_nl = ~ or_tmp_529;
  assign rec_quad_normal_x_not_nl = ~ or_tmp_529;
  assign nl_quadInters_run_if_2_acc_nl = conv_s2u_34_35(ac_math_ac_abs_58_58_xabs_acc_itm_57_24)
      + 35'b11111111111111111111111111111111001;
  assign quadInters_run_if_2_acc_nl = nl_quadInters_run_if_2_acc_nl[34:0];
  assign nl_quadInters_denom_dot_run_acc_2_nl = (quadInters_denom_dot_run_mul_1_cmp_z_oreg[57:0])
      + quadInters_denom_dot_run_mul_2_cmp_z_oreg;
  assign quadInters_denom_dot_run_acc_2_nl = nl_quadInters_denom_dot_run_acc_2_nl[57:0];
  assign ac_math_ac_abs_58_58_xabs_xor_nl = (signext_58_1(quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0[57]))
      ^ quadInters_denom_dot_run_ac_fixed_cctor_sva_mx2w0;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_30_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_61_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1[34]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl
      = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_32_sva_1[33:0])
      , div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_2_itm_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_30_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_61_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_32_acc_1_nl[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_62_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_mx1w0,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1[33]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl
      = ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_1_acc_1_psp_sva_1
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_mx0_33_32[0])})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_62_nl)});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_2_acc_1_nl[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_4_nl
      = (~ quadInters_run_if_2_slc_quadInters_run_if_2_acc_34_svs) & (fsm_output[5]);
  assign setfacenorm_dot_run_and_1_nl = (~ quadInters_run_lor_3_lpi_2_dfm) & (fsm_output[5]);
  assign nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl
      = conv_u2u_33_34(~ quadInters_run_rounded_denom_lpi_2_dfm_mx0_32_0) + 34'b0000000000000000000000000000000001;
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl
      = nl_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qif_acc_nl[33:0];
  assign quadInters_cross_v_run_mul_6_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg , (add_run_ac_fixed_cctor_2_74_43_sva[8:0])
      , (mult_run_asn_2_itm_1_74_30[12:0])})) * $signed((quads_crt_sva_7_110_0[83:72])));
  assign quadInters_cross_v_run_mux_2_nl = MUX_v_60_2_2((signext_60_57(quadInters_cross_v_run_mul_6_nl)),
      setfacenorm_dot_run_acc_2_itm, fsm_output[2]);
  assign quadInters_cross_v_run_or_1_nl = (~ (fsm_output[2])) | (fsm_output[4]);
  assign quadInters_cross_v_run_mul_7_nl = conv_s2u_57_57($signed(({reg_quadInters_sub_run_ac_fixed_cctor_44_22_reg
      , reg_quadInters_sub_run_ac_fixed_cctor_44_22_1_reg , (add_run_ac_fixed_cctor_74_43_sva[8:0])
      , quadInters_at_run_mult_result_x_74_30_sva_12_0})) * $signed((quads_crt_sva_7_110_0[107:96])));
  assign quadInters_cross_v_run_mux_3_nl = MUX_v_60_2_2((signext_60_57(~ (quadInters_cross_v_run_mul_7_nl))),
      quadInters_denom_dot_run_mul_1_cmp_z_oreg, fsm_output[2]);
  assign nl_acc_nl = ({(quadInters_cross_v_run_mux_2_nl) , (quadInters_cross_v_run_or_1_nl)})
      + ({(quadInters_cross_v_run_mux_3_nl) , 1'b1});
  assign acc_nl = nl_acc_nl[60:0];
  assign z_out = readslicef_61_60_1((acc_nl));
  assign for_for_and_2_nl = MUX_v_15_2_2(15'b000000000000000, (reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1[19:5]),
      (fsm_output[3]));
  assign for_mux_25_nl = MUX_v_5_2_2(for_i_5_0_sva_4_0, (reg_ac_math_ac_abs_21_21_2_xabs_xor_ftd_1[4:0]),
      fsm_output[3]);
  assign for_or_11_nl = (reg_quadInters_sub_run_ac_fixed_cctor_2_44_22_1_reg[20])
      | (fsm_output[2]);
  assign nl_z_out_1 = conv_u2u_20_21({(for_for_and_2_nl) , (for_mux_25_nl)}) + conv_u2u_1_21(for_or_11_nl);
  assign z_out_1 = nl_z_out_1[20:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_21_nl
      = (fsm_output[2]) | (fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1[32:0]),
      (z_out_5[32:0]), div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_21_nl);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_131_nl
      = MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_50_lpi_2_dfm_mx0[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_40_lpi_2_dfm_mx0[0]),
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_82_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_35_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_83_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (z_out_5[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_84_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (z_out_5[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_132_nl
      = MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_82_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_83_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_84_nl),
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_133_nl
      = MUX1HOT_v_33_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_68_lpi_2_dfm_mx0[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx1[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx3[33:1]),
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4])});
  assign nl_z_out_2 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_131_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_132_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_133_nl)});
  assign z_out_2 = nl_z_out_2[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_85_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1[33])
      & (~ (fsm_output[4]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_123_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1[32:0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1[32:0]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_124_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_61_lpi_2_dfm_mx0[0]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_86_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_126_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_12_sva_1[34]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_87_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_29_psp_sva_mx0w1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_125_nl
      = MUX_v_35_2_2(({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_86_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_126_nl)}),
      (signext_35_34({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_87_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_37_lpi_2_dfm_mx2[33:1])})),
      fsm_output[4]);
  assign nl_z_out_3 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_85_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_123_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_124_nl)})
      + (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_125_nl);
  assign z_out_3 = nl_z_out_3[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_127_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[32:0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1[32:0]),
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_128_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_45_lpi_2_dfm_mx0[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_35_lpi_2_dfm_mx0[0]),
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_88_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_13_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_89_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_3_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_129_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_88_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_89_nl),
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_130_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_46_lpi_2_dfm_mx0[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_mx2[33:1]),
      fsm_output[3]);
  assign nl_z_out_4 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_127_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_128_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_129_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_130_nl)});
  assign z_out_4 = nl_z_out_4[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_131_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1[32:0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1[32:0]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_132_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_49_lpi_2_dfm_mx0[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_39_lpi_2_dfm_mx0[0]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_90_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_17_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_91_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_7_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_133_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_90_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_91_nl),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_134_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_50_lpi_2_dfm_mx0[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_40_lpi_2_dfm_mx0[33:1]),
      fsm_output[4]);
  assign nl_z_out_5 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_131_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_132_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_133_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_134_nl)});
  assign z_out_5 = nl_z_out_5[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_135_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[32:0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[32:0]),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_136_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_59_lpi_2_dfm_mx0[0]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_65_lpi_2_dfm_mx0[0]),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_92_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_27_psp_sva_mx0w2[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_93_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_33_psp_sva_1[33]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_137_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_92_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_93_nl),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_138_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_60_lpi_2_dfm_mx0[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_66_lpi_2_dfm_mx0[33:1]),
      fsm_output[5]);
  assign nl_z_out_6 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_135_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_136_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_137_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_138_nl)});
  assign z_out_6 = nl_z_out_6[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_94_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_3[33])
      & (~ div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_sva_33);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_95_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_41_psp_ftd);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_139_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_94_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_95_nl),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_140_nl
      = MUX_v_33_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_52_lpi_2_dfm_mx0[33:1]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_42_lpi_2_dfm_mx0[33:1]),
      fsm_output[5]);
  assign nl_z_out_7 = ({reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_acc_19_psp_1_cse
      , reg_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_qr_33_0_36_lpi_2_dfm_ftd_1})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_139_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_140_nl)});
  assign z_out_7 = nl_z_out_7[33:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_14_nl
      = MUX_v_34_2_2((z_out_13[33:0]), (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1[33:0]),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_134_nl
      = MUX1HOT_s_1_3_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[17]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[12]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[7]),
      {(fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_96_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_13[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_97_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_15_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_96_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_97_nl),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_22_nl
      = ((z_out_13[34]) & (fsm_output[3])) | ((z_out_13[34]) & (fsm_output[4])) |
      ((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_27_sva_1[34])
      & (fsm_output[5]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_16_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_22_nl);
  assign nl_z_out_8 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_14_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_134_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_15_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_16_nl)});
  assign z_out_8 = nl_z_out_8[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_141_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[20]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[10]),
      fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_23_nl
      = ((z_out_10[34]) & (~ (fsm_output[5]))) | ((z_out_10[34]) & (fsm_output[5]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_142_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_23_nl);
  assign nl_z_out_9 = ({(z_out_10[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_141_nl)})
      + ({div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_12_cse
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_142_nl)});
  assign z_out_9 = nl_z_out_9[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_135_nl
      = MUX1HOT_s_1_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_6_itm_1,
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[21]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[16]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[11]),
      {(fsm_output[2]) , (fsm_output[3]) , (fsm_output[4]) , (fsm_output[5])});
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_98_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_99_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_98_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_99_nl),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_m1c);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_24_nl
      = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl
      = (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34]))
      & (fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[34])
      & (fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_136_nl
      = MUX1HOT_v_34_3_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_33_itm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      {(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_24_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_47_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_48_nl)});
  assign nl_z_out_10 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_13_sva[33:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_135_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_17_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_136_nl)});
  assign z_out_10 = nl_z_out_10[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_143_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22[3]),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_35_operator_35_true_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_R_34_1_itm,
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_100_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_12[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_101_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (z_out_12[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_144_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_100_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_101_nl),
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_145_nl
      = MUX_v_34_4_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      {(fsm_output[3]) , (z_out_12[34])});
  assign nl_z_out_11 = ({(z_out_12[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_143_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_144_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_145_nl)});
  assign z_out_11 = nl_z_out_11[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_146_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_26_22[4]),
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_N_slc_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_1_itm_1,
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_102_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_103_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_147_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_102_nl),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_103_nl),
      fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_49_nl
      = (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34]))
      & (fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_50_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[34])
      & (fsm_output[3]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_2_nl
      = MUX1HOT_v_34_3_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_13_itm,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_2,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_2,
      {(~ (fsm_output[3])) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_49_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_50_nl)});
  assign nl_z_out_12 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_3_sva[33:0])
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_146_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_147_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux1h_2_nl)});
  assign z_out_12 = nl_z_out_12[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_148_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[18]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[13]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_104_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (z_out_14[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_25_nl
      = ((z_out_14[34]) & (~ (fsm_output[4]))) | ((z_out_14[34]) & (fsm_output[4]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_149_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_25_nl);
  assign nl_z_out_13 = ({(z_out_14[33:0]) , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_148_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_104_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_149_nl)});
  assign z_out_13 = nl_z_out_13[34:0];
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_150_nl
      = MUX_v_34_2_2((z_out_9[33:0]), (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1[33:0]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_151_nl
      = MUX_s_1_2_2((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[19]),
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uN_qr_lpi_2_dfm_1_21_0[14]),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_105_nl
      = (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1[33])
      & (~ (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1[34]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_152_nl
      = MUX_s_1_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_13_cse,
      (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_and_105_nl),
      fsm_output[4]);
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_26_nl
      = ((z_out_9[34]) & (~ (fsm_output[4]))) | ((div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_ac_int_cctor_20_sva_1[34])
      & (fsm_output[4]));
  assign div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_153_nl
      = MUX_v_34_2_2(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_neg_D_acc_psp_sva_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_uD_qr_lpi_2_dfm_1,
      div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_or_26_nl);
  assign nl_z_out_14 = ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_150_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_151_nl)})
      + ({(div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_152_nl)
      , (div_34_14_AC_TRN_AC_WRAP_34_11_AC_TRN_AC_WRAP_60_17_AC_TRN_AC_WRAP_1_for_mux_153_nl)});
  assign z_out_14 = nl_z_out_14[34:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_3_2;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [2:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | ( input_1 & {26{sel[1]}});
    result = result | ( input_2 & {26{sel[2]}});
    MUX1HOT_v_26_3_2 = result;
  end
  endfunction


  function automatic [25:0] MUX1HOT_v_26_4_2;
    input [25:0] input_3;
    input [25:0] input_2;
    input [25:0] input_1;
    input [25:0] input_0;
    input [3:0] sel;
    reg [25:0] result;
  begin
    result = input_0 & {26{sel[0]}};
    result = result | ( input_1 & {26{sel[1]}});
    result = result | ( input_2 & {26{sel[2]}});
    result = result | ( input_3 & {26{sel[3]}});
    MUX1HOT_v_26_4_2 = result;
  end
  endfunction


  function automatic [32:0] MUX1HOT_v_33_3_2;
    input [32:0] input_2;
    input [32:0] input_1;
    input [32:0] input_0;
    input [2:0] sel;
    reg [32:0] result;
  begin
    result = input_0 & {33{sel[0]}};
    result = result | ( input_1 & {33{sel[1]}});
    result = result | ( input_2 & {33{sel[2]}});
    MUX1HOT_v_33_3_2 = result;
  end
  endfunction


  function automatic [33:0] MUX1HOT_v_34_3_2;
    input [33:0] input_2;
    input [33:0] input_1;
    input [33:0] input_0;
    input [2:0] sel;
    reg [33:0] result;
  begin
    result = input_0 & {34{sel[0]}};
    result = result | ( input_1 & {34{sel[1]}});
    result = result | ( input_2 & {34{sel[2]}});
    MUX1HOT_v_34_3_2 = result;
  end
  endfunction


  function automatic [33:0] MUX1HOT_v_34_4_2;
    input [33:0] input_3;
    input [33:0] input_2;
    input [33:0] input_1;
    input [33:0] input_0;
    input [3:0] sel;
    reg [33:0] result;
  begin
    result = input_0 & {34{sel[0]}};
    result = result | ( input_1 & {34{sel[1]}});
    result = result | ( input_2 & {34{sel[2]}});
    result = result | ( input_3 & {34{sel[3]}});
    MUX1HOT_v_34_4_2 = result;
  end
  endfunction


  function automatic [34:0] MUX1HOT_v_35_3_2;
    input [34:0] input_2;
    input [34:0] input_1;
    input [34:0] input_0;
    input [2:0] sel;
    reg [34:0] result;
  begin
    result = input_0 & {35{sel[0]}};
    result = result | ( input_1 & {35{sel[1]}});
    result = result | ( input_2 & {35{sel[2]}});
    MUX1HOT_v_35_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input [0:0] sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction


  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function automatic [24:0] MUX_v_25_2_2;
    input [24:0] input_0;
    input [24:0] input_1;
    input [0:0] sel;
    reg [24:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_25_2_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_2_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input [0:0] sel;
    reg [25:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_26_2_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_2_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input [0:0] sel;
    reg [26:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_27_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [32:0] MUX_v_33_2_2;
    input [32:0] input_0;
    input [32:0] input_1;
    input [0:0] sel;
    reg [32:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_33_2_2 = result;
  end
  endfunction


  function automatic [33:0] MUX_v_34_2_2;
    input [33:0] input_0;
    input [33:0] input_1;
    input [0:0] sel;
    reg [33:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_34_2_2 = result;
  end
  endfunction


  function automatic [33:0] MUX_v_34_4_2;
    input [33:0] input_0;
    input [33:0] input_1;
    input [33:0] input_2;
    input [33:0] input_3;
    input [1:0] sel;
    reg [33:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      2'b10 : begin
        result = input_2;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_34_4_2 = result;
  end
  endfunction


  function automatic [34:0] MUX_v_35_2_2;
    input [34:0] input_0;
    input [34:0] input_1;
    input [0:0] sel;
    reg [34:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_35_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [55:0] MUX_v_56_2_2;
    input [55:0] input_0;
    input [55:0] input_1;
    input [0:0] sel;
    reg [55:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_56_2_2 = result;
  end
  endfunction


  function automatic [57:0] MUX_v_58_2_2;
    input [57:0] input_0;
    input [57:0] input_1;
    input [0:0] sel;
    reg [57:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_58_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [59:0] MUX_v_60_2_2;
    input [59:0] input_0;
    input [59:0] input_1;
    input [0:0] sel;
    reg [59:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_60_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_22_1_21;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 21;
    readslicef_22_1_21 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_28_1_27;
    input [27:0] vector;
    reg [27:0] tmp;
  begin
    tmp = vector >> 27;
    readslicef_28_1_27 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_35_1_34;
    input [34:0] vector;
    reg [34:0] tmp;
  begin
    tmp = vector >> 34;
    readslicef_35_1_34 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_39_1_38;
    input [38:0] vector;
    reg [38:0] tmp;
  begin
    tmp = vector >> 38;
    readslicef_39_1_38 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_48_1_47;
    input [47:0] vector;
    reg [47:0] tmp;
  begin
    tmp = vector >> 47;
    readslicef_48_1_47 = tmp[0:0];
  end
  endfunction


  function automatic [33:0] readslicef_48_34_14;
    input [47:0] vector;
    reg [47:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_48_34_14 = tmp[33:0];
  end
  endfunction


  function automatic [55:0] readslicef_57_56_1;
    input [56:0] vector;
    reg [56:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_57_56_1 = tmp[55:0];
  end
  endfunction


  function automatic [33:0] readslicef_58_34_24;
    input [57:0] vector;
    reg [57:0] tmp;
  begin
    tmp = vector >> 24;
    readslicef_58_34_24 = tmp[33:0];
  end
  endfunction


  function automatic [0:0] readslicef_60_1_59;
    input [59:0] vector;
    reg [59:0] tmp;
  begin
    tmp = vector >> 59;
    readslicef_60_1_59 = tmp[0:0];
  end
  endfunction


  function automatic [46:0] readslicef_60_47_13;
    input [59:0] vector;
    reg [59:0] tmp;
  begin
    tmp = vector >> 13;
    readslicef_60_47_13 = tmp[46:0];
  end
  endfunction


  function automatic [59:0] readslicef_61_60_1;
    input [60:0] vector;
    reg [60:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_61_60_1 = tmp[59:0];
  end
  endfunction


  function automatic [37:0] readslicef_62_38_24;
    input [61:0] vector;
    reg [61:0] tmp;
  begin
    tmp = vector >> 24;
    readslicef_62_38_24 = tmp[37:0];
  end
  endfunction


  function automatic [19:0] signext_20_1;
    input [0:0] vector;
  begin
    signext_20_1= {{19{vector[0]}}, vector};
  end
  endfunction


  function automatic [24:0] signext_25_21;
    input [20:0] vector;
  begin
    signext_25_21= {{4{vector[20]}}, vector};
  end
  endfunction


  function automatic [34:0] signext_35_34;
    input [33:0] vector;
  begin
    signext_35_34= {{1{vector[33]}}, vector};
  end
  endfunction


  function automatic [55:0] signext_56_26;
    input [25:0] vector;
  begin
    signext_56_26= {{30{vector[25]}}, vector};
  end
  endfunction


  function automatic [57:0] signext_58_1;
    input [0:0] vector;
  begin
    signext_58_1= {{57{vector[0]}}, vector};
  end
  endfunction


  function automatic [59:0] signext_60_57;
    input [56:0] vector;
  begin
    signext_60_57= {{3{vector[56]}}, vector};
  end
  endfunction


  function automatic [33:0] conv_s2s_31_34 ;
    input [30:0]  vector ;
  begin
    conv_s2s_31_34 = {{3{vector[30]}}, vector};
  end
  endfunction


  function automatic [38:0] conv_s2s_38_39 ;
    input [37:0]  vector ;
  begin
    conv_s2s_38_39 = {vector[37], vector};
  end
  endfunction


  function automatic [47:0] conv_s2s_47_48 ;
    input [46:0]  vector ;
  begin
    conv_s2s_47_48 = {vector[46], vector};
  end
  endfunction


  function automatic [22:0] conv_s2u_12_23 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_23 = {{11{vector[11]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [31:0] conv_s2u_21_32 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_32 = {{11{vector[20]}}, vector};
  end
  endfunction


  function automatic [27:0] conv_s2u_27_28 ;
    input [26:0]  vector ;
  begin
    conv_s2u_27_28 = {vector[26], vector};
  end
  endfunction


  function automatic [34:0] conv_s2u_34_35 ;
    input [33:0]  vector ;
  begin
    conv_s2u_34_35 = {vector[33], vector};
  end
  endfunction


  function automatic [47:0] conv_s2u_47_48 ;
    input [46:0]  vector ;
  begin
    conv_s2u_47_48 = {vector[46], vector};
  end
  endfunction


  function automatic [56:0] conv_s2u_57_57 ;
    input [56:0]  vector ;
  begin
    conv_s2u_57_57 = vector;
  end
  endfunction


  function automatic [20:0] conv_u2s_1_21 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_21 = {{20{1'b0}}, vector};
  end
  endfunction


  function automatic [33:0] conv_u2s_1_34 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_34 = {{33{1'b0}}, vector};
  end
  endfunction


  function automatic [59:0] conv_u2s_1_60 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_60 = {{59{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [20:0] conv_u2s_20_21 ;
    input [19:0]  vector ;
  begin
    conv_u2s_20_21 =  {1'b0, vector};
  end
  endfunction


  function automatic [34:0] conv_u2s_34_35 ;
    input [33:0]  vector ;
  begin
    conv_u2s_34_35 =  {1'b0, vector};
  end
  endfunction


  function automatic [20:0] conv_u2u_1_21 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_21 = {{20{1'b0}}, vector};
  end
  endfunction


  function automatic [57:0] conv_u2u_1_58 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_58 = {{57{1'b0}}, vector};
  end
  endfunction


  function automatic [20:0] conv_u2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_u2u_20_21 = {1'b0, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit_hit
// ------------------------------------------------------------------


module WorldHit_hit (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld,
      attenuation_chan_in_rsc_rdy, accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld,
      accumalated_color_chan_in_rsc_rdy, quad_hit_anything_outone_rsc_dat, quad_hit_anything_outone_rsc_vld,
      quad_hit_anything_outone_rsc_rdy, quad_hit_anything_outtwo_rsc_dat, quad_hit_anything_outtwo_rsc_vld,
      quad_hit_anything_outtwo_rsc_rdy, rec_quad_outone_rsc_dat, rec_quad_outone_rsc_vld,
      rec_quad_outone_rsc_rdy, rec_quad_outtwo_rsc_dat, rec_quad_outtwo_rsc_vld,
      rec_quad_outtwo_rsc_rdy, closest_so_far_outone_rsc_dat, closest_so_far_outone_rsc_vld,
      closest_so_far_outone_rsc_rdy, closest_so_far_outtwo_rsc_dat, closest_so_far_outtwo_rsc_vld,
      closest_so_far_outtwo_rsc_rdy, attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld,
      attenuation_chan_out_rsc_rdy, accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld,
      accumalated_color_out_rsc_rdy, hit_out_rsc_dat, hit_out_rsc_vld, hit_out_rsc_rdy,
      ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, isHit_rsc_dat, isHit_rsc_vld,
      isHit_rsc_rdy, else_mul_cmp_a, else_mul_cmp_b, else_mul_cmp_z
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input quad_hit_anything_outone_rsc_dat;
  input quad_hit_anything_outone_rsc_vld;
  output quad_hit_anything_outone_rsc_rdy;
  input quad_hit_anything_outtwo_rsc_dat;
  input quad_hit_anything_outtwo_rsc_vld;
  output quad_hit_anything_outtwo_rsc_rdy;
  input [225:0] rec_quad_outone_rsc_dat;
  input rec_quad_outone_rsc_vld;
  output rec_quad_outone_rsc_rdy;
  input [225:0] rec_quad_outtwo_rsc_dat;
  input rec_quad_outtwo_rsc_vld;
  output rec_quad_outtwo_rsc_rdy;
  input [46:0] closest_so_far_outone_rsc_dat;
  input closest_so_far_outone_rsc_vld;
  output closest_so_far_outone_rsc_rdy;
  input [46:0] closest_so_far_outtwo_rsc_dat;
  input closest_so_far_outtwo_rsc_vld;
  output closest_so_far_outtwo_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [225:0] hit_out_rsc_dat;
  output hit_out_rsc_vld;
  input hit_out_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  output isHit_rsc_dat;
  output isHit_rsc_vld;
  input isHit_rsc_rdy;
  output [26:0] else_mul_cmp_a;
  reg [26:0] else_mul_cmp_a;
  output [26:0] else_mul_cmp_b;
  reg [26:0] else_mul_cmp_b;
  input [48:0] else_mul_cmp_z;


  // Interconnect Declarations
  wire hit_wen;
  wire ray_in_rsci_wen_comp;
  wire [164:0] ray_in_rsci_idat_mxwt;
  wire params_in_rsci_wen_comp;
  wire [80:0] params_in_rsci_idat_mxwt;
  wire attenuation_chan_in_rsci_wen_comp;
  wire [80:0] attenuation_chan_in_rsci_idat_mxwt;
  wire accumalated_color_chan_in_rsci_wen_comp;
  wire [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  wire quad_hit_anything_outone_rsci_wen_comp;
  wire quad_hit_anything_outone_rsci_idat_mxwt;
  wire quad_hit_anything_outtwo_rsci_wen_comp;
  wire quad_hit_anything_outtwo_rsci_idat_mxwt;
  wire rec_quad_outone_rsci_wen_comp;
  wire [225:0] rec_quad_outone_rsci_idat_mxwt;
  wire rec_quad_outtwo_rsci_wen_comp;
  wire [225:0] rec_quad_outtwo_rsci_idat_mxwt;
  wire closest_so_far_outone_rsci_wen_comp;
  wire [46:0] closest_so_far_outone_rsci_idat_mxwt;
  wire closest_so_far_outtwo_rsci_wen_comp;
  wire [46:0] closest_so_far_outtwo_rsci_idat_mxwt;
  wire attenuation_chan_out_rsci_wen_comp;
  reg [80:0] attenuation_chan_out_rsci_idat;
  wire accumalated_color_out_rsci_wen_comp;
  wire hit_out_rsci_wen_comp;
  wire ray_out_rsci_wen_comp;
  wire isHit_rsci_wen_comp;
  wire [26:0] else_mul_cmp_z_oreg;
  reg [26:0] accumalated_color_out_rsci_idat_80_54;
  reg [26:0] accumalated_color_out_rsci_idat_53_27;
  reg [26:0] accumalated_color_out_rsci_idat_26_0;
  reg [26:0] hit_out_rsci_idat_225_199;
  reg [26:0] hit_out_rsci_idat_198_172;
  reg [26:0] hit_out_rsci_idat_171_145;
  reg [2:0] hit_out_rsci_idat_144_142;
  reg hit_out_rsci_idat_141;
  reg [25:0] hit_out_rsci_idat_140_115;
  reg [25:0] hit_out_rsci_idat_114_89;
  reg [25:0] hit_out_rsci_idat_88_63;
  reg [20:0] hit_out_rsci_idat_62_42;
  reg [20:0] hit_out_rsci_idat_41_21;
  reg [20:0] hit_out_rsci_idat_20_0;
  reg [164:0] ray_out_rsci_idat_164_0;
  wire [6:0] fsm_output;
  wire and_dcpl;
  wire ray_out_and_cse;
  wire accumalated_color_out_and_cse;
  reg reg_isHit_rsci_ivld_hit_psct_cse;
  reg reg_accumalated_color_out_rsci_ivld_hit_psct_cse;
  reg reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse;
  wire [26:0] z_out;
  wire [27:0] nl_z_out;
  reg [80:0] accumalated_color_chan_in_crt_sva;
  reg if_slc_47_svs;
  reg [26:0] mux_12_itm;
  reg [26:0] mux_11_itm;
  wire or_mdf_sva_mx0w0;
  reg reg_isHit_rsci_idat_cse;
  reg [26:0] attenuation_chan_in_crt_sva_80_54;
  reg [26:0] attenuation_chan_in_crt_sva_53_27;
  reg [26:0] params_in_crt_sva_91_65;
  reg [26:0] params_in_crt_sva_64_38;
  wire and_94_cse;
  wire if_acc_itm_47;

  wire[20:0] if_mux_nl;
  wire[20:0] if_mux_1_nl;
  wire[20:0] if_mux_2_nl;
  wire[25:0] if_mux_3_nl;
  wire[25:0] if_mux_4_nl;
  wire[25:0] if_mux_5_nl;
  wire[0:0] if_mux_6_nl;
  wire[0:0] if_if_mux_1_nl;
  wire[2:0] if_mux_7_nl;
  wire[26:0] if_mux_8_nl;
  wire[26:0] if_mux_9_nl;
  wire[26:0] if_mux_10_nl;
  wire[0:0] and_45_nl;
  wire[0:0] and_82_nl;
  wire[47:0] if_acc_nl;
  wire[48:0] nl_if_acc_nl;
  wire[26:0] else_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [80:0] nl_WorldHit_hit_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat;
  assign nl_WorldHit_hit_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat
      = {accumalated_color_out_rsci_idat_80_54 , accumalated_color_out_rsci_idat_53_27
      , accumalated_color_out_rsci_idat_26_0};
  wire [225:0] nl_WorldHit_hit_hit_out_rsci_inst_hit_out_rsci_idat;
  assign nl_WorldHit_hit_hit_out_rsci_inst_hit_out_rsci_idat = {hit_out_rsci_idat_225_199
      , hit_out_rsci_idat_198_172 , hit_out_rsci_idat_171_145 , hit_out_rsci_idat_144_142
      , hit_out_rsci_idat_141 , hit_out_rsci_idat_140_115 , hit_out_rsci_idat_114_89
      , hit_out_rsci_idat_88_63 , hit_out_rsci_idat_62_42 , hit_out_rsci_idat_41_21
      , hit_out_rsci_idat_20_0};
  wire [165:0] nl_WorldHit_hit_ray_out_rsci_inst_ray_out_rsci_idat;
  assign nl_WorldHit_hit_ray_out_rsci_inst_ray_out_rsci_idat = {1'b0 , ray_out_rsci_idat_164_0};
  WorldHit_hit_ray_in_rsci WorldHit_hit_ray_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .hit_wen(hit_wen),
      .ray_in_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt)
    );
  WorldHit_hit_params_in_rsci WorldHit_hit_params_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .hit_wen(hit_wen),
      .params_in_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt)
    );
  WorldHit_hit_attenuation_chan_in_rsci WorldHit_hit_attenuation_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .hit_wen(hit_wen),
      .attenuation_chan_in_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt)
    );
  WorldHit_hit_accumalated_color_chan_in_rsci WorldHit_hit_accumalated_color_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .hit_wen(hit_wen),
      .accumalated_color_chan_in_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt)
    );
  WorldHit_hit_quad_hit_anything_outone_rsci WorldHit_hit_quad_hit_anything_outone_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_outone_rsc_dat(quad_hit_anything_outone_rsc_dat),
      .quad_hit_anything_outone_rsc_vld(quad_hit_anything_outone_rsc_vld),
      .quad_hit_anything_outone_rsc_rdy(quad_hit_anything_outone_rsc_rdy),
      .hit_wen(hit_wen),
      .quad_hit_anything_outone_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .quad_hit_anything_outone_rsci_wen_comp(quad_hit_anything_outone_rsci_wen_comp),
      .quad_hit_anything_outone_rsci_idat_mxwt(quad_hit_anything_outone_rsci_idat_mxwt)
    );
  WorldHit_hit_quad_hit_anything_outtwo_rsci WorldHit_hit_quad_hit_anything_outtwo_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .quad_hit_anything_outtwo_rsc_dat(quad_hit_anything_outtwo_rsc_dat),
      .quad_hit_anything_outtwo_rsc_vld(quad_hit_anything_outtwo_rsc_vld),
      .quad_hit_anything_outtwo_rsc_rdy(quad_hit_anything_outtwo_rsc_rdy),
      .hit_wen(hit_wen),
      .quad_hit_anything_outtwo_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .quad_hit_anything_outtwo_rsci_wen_comp(quad_hit_anything_outtwo_rsci_wen_comp),
      .quad_hit_anything_outtwo_rsci_idat_mxwt(quad_hit_anything_outtwo_rsci_idat_mxwt)
    );
  WorldHit_hit_rec_quad_outone_rsci WorldHit_hit_rec_quad_outone_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_outone_rsc_dat(rec_quad_outone_rsc_dat),
      .rec_quad_outone_rsc_vld(rec_quad_outone_rsc_vld),
      .rec_quad_outone_rsc_rdy(rec_quad_outone_rsc_rdy),
      .hit_wen(hit_wen),
      .rec_quad_outone_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .rec_quad_outone_rsci_wen_comp(rec_quad_outone_rsci_wen_comp),
      .rec_quad_outone_rsci_idat_mxwt(rec_quad_outone_rsci_idat_mxwt)
    );
  WorldHit_hit_rec_quad_outtwo_rsci WorldHit_hit_rec_quad_outtwo_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rec_quad_outtwo_rsc_dat(rec_quad_outtwo_rsc_dat),
      .rec_quad_outtwo_rsc_vld(rec_quad_outtwo_rsc_vld),
      .rec_quad_outtwo_rsc_rdy(rec_quad_outtwo_rsc_rdy),
      .hit_wen(hit_wen),
      .rec_quad_outtwo_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .rec_quad_outtwo_rsci_wen_comp(rec_quad_outtwo_rsci_wen_comp),
      .rec_quad_outtwo_rsci_idat_mxwt(rec_quad_outtwo_rsci_idat_mxwt)
    );
  WorldHit_hit_closest_so_far_outone_rsci WorldHit_hit_closest_so_far_outone_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_outone_rsc_dat(closest_so_far_outone_rsc_dat),
      .closest_so_far_outone_rsc_vld(closest_so_far_outone_rsc_vld),
      .closest_so_far_outone_rsc_rdy(closest_so_far_outone_rsc_rdy),
      .hit_wen(hit_wen),
      .closest_so_far_outone_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .closest_so_far_outone_rsci_wen_comp(closest_so_far_outone_rsci_wen_comp),
      .closest_so_far_outone_rsci_idat_mxwt(closest_so_far_outone_rsci_idat_mxwt)
    );
  WorldHit_hit_closest_so_far_outtwo_rsci WorldHit_hit_closest_so_far_outtwo_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .closest_so_far_outtwo_rsc_dat(closest_so_far_outtwo_rsc_dat),
      .closest_so_far_outtwo_rsc_vld(closest_so_far_outtwo_rsc_vld),
      .closest_so_far_outtwo_rsc_rdy(closest_so_far_outtwo_rsc_rdy),
      .hit_wen(hit_wen),
      .closest_so_far_outtwo_rsci_oswt(reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse),
      .closest_so_far_outtwo_rsci_wen_comp(closest_so_far_outtwo_rsci_wen_comp),
      .closest_so_far_outtwo_rsci_idat_mxwt(closest_so_far_outtwo_rsci_idat_mxwt)
    );
  WorldHit_hit_attenuation_chan_out_rsci WorldHit_hit_attenuation_chan_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .hit_wen(hit_wen),
      .attenuation_chan_out_rsci_oswt(reg_isHit_rsci_ivld_hit_psct_cse),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_idat(attenuation_chan_out_rsci_idat)
    );
  WorldHit_hit_accumalated_color_out_rsci WorldHit_hit_accumalated_color_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .hit_wen(hit_wen),
      .accumalated_color_out_rsci_oswt(reg_accumalated_color_out_rsci_ivld_hit_psct_cse),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_idat(nl_WorldHit_hit_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat[80:0])
    );
  WorldHit_hit_hit_out_rsci WorldHit_hit_hit_out_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .hit_out_rsc_dat(hit_out_rsc_dat),
      .hit_out_rsc_vld(hit_out_rsc_vld),
      .hit_out_rsc_rdy(hit_out_rsc_rdy),
      .hit_wen(hit_wen),
      .hit_out_rsci_oswt(reg_isHit_rsci_ivld_hit_psct_cse),
      .hit_out_rsci_wen_comp(hit_out_rsci_wen_comp),
      .hit_out_rsci_idat(nl_WorldHit_hit_hit_out_rsci_inst_hit_out_rsci_idat[225:0])
    );
  WorldHit_hit_ray_out_rsci WorldHit_hit_ray_out_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .hit_wen(hit_wen),
      .ray_out_rsci_oswt(reg_isHit_rsci_ivld_hit_psct_cse),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_idat(nl_WorldHit_hit_ray_out_rsci_inst_ray_out_rsci_idat[165:0])
    );
  WorldHit_hit_isHit_rsci WorldHit_hit_isHit_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .isHit_rsc_dat(isHit_rsc_dat),
      .isHit_rsc_vld(isHit_rsc_vld),
      .isHit_rsc_rdy(isHit_rsc_rdy),
      .hit_wen(hit_wen),
      .isHit_rsci_oswt(reg_isHit_rsci_ivld_hit_psct_cse),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp),
      .isHit_rsci_idat(reg_isHit_rsci_idat_cse)
    );
  WorldHit_hit_wait_dp WorldHit_hit_wait_dp_inst (
      .clk(clk),
      .arst_n(arst_n),
      .else_mul_cmp_z(else_mul_cmp_z),
      .hit_wen(hit_wen),
      .else_mul_cmp_z_oreg(else_mul_cmp_z_oreg)
    );
  WorldHit_hit_staller WorldHit_hit_staller_inst (
      .hit_wen(hit_wen),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .quad_hit_anything_outone_rsci_wen_comp(quad_hit_anything_outone_rsci_wen_comp),
      .quad_hit_anything_outtwo_rsci_wen_comp(quad_hit_anything_outtwo_rsci_wen_comp),
      .rec_quad_outone_rsci_wen_comp(rec_quad_outone_rsci_wen_comp),
      .rec_quad_outtwo_rsci_wen_comp(rec_quad_outtwo_rsci_wen_comp),
      .closest_so_far_outone_rsci_wen_comp(closest_so_far_outone_rsci_wen_comp),
      .closest_so_far_outtwo_rsci_wen_comp(closest_so_far_outtwo_rsci_wen_comp),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .hit_out_rsci_wen_comp(hit_out_rsci_wen_comp),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp)
    );
  WorldHit_hit_hit_fsm WorldHit_hit_hit_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .hit_wen(hit_wen),
      .fsm_output(fsm_output)
    );
  assign ray_out_and_cse = hit_wen & (fsm_output[1]);
  assign accumalated_color_out_and_cse = hit_wen & (fsm_output[5]);
  assign and_94_cse = (~ (fsm_output[2])) & hit_wen;
  assign or_mdf_sva_mx0w0 = quad_hit_anything_outone_rsci_idat_mxwt | quad_hit_anything_outtwo_rsci_idat_mxwt;
  assign nl_if_acc_nl = conv_s2u_47_48(closest_so_far_outone_rsci_idat_mxwt) - conv_s2u_47_48(closest_so_far_outtwo_rsci_idat_mxwt);
  assign if_acc_nl = nl_if_acc_nl[47:0];
  assign if_acc_itm_47 = readslicef_48_1_47((if_acc_nl));
  assign and_dcpl = ~(quad_hit_anything_outtwo_rsci_idat_mxwt | quad_hit_anything_outone_rsci_idat_mxwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_rsci_idat_164_0 <= 165'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      hit_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      hit_out_rsci_idat_41_21 <= 21'b000000000000000000000;
      hit_out_rsci_idat_62_42 <= 21'b000000000000000000000;
      hit_out_rsci_idat_88_63 <= 26'b00000000000000000000000000;
      hit_out_rsci_idat_114_89 <= 26'b00000000000000000000000000;
      hit_out_rsci_idat_140_115 <= 26'b00000000000000000000000000;
      hit_out_rsci_idat_141 <= 1'b0;
      hit_out_rsci_idat_144_142 <= 3'b000;
      hit_out_rsci_idat_171_145 <= 27'b000000000000000000000000000;
      hit_out_rsci_idat_198_172 <= 27'b000000000000000000000000000;
      hit_out_rsci_idat_225_199 <= 27'b000000000000000000000000000;
      reg_isHit_rsci_idat_cse <= 1'b0;
      attenuation_chan_out_rsci_idat <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      accumalated_color_chan_in_crt_sva <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ray_out_and_cse ) begin
      ray_out_rsci_idat_164_0 <= ray_in_rsci_idat_mxwt;
      hit_out_rsci_idat_20_0 <= MUX_v_21_2_2(21'b000000000000000000000, (if_mux_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_41_21 <= MUX_v_21_2_2(21'b000000000000000000000, (if_mux_1_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_62_42 <= MUX_v_21_2_2(21'b000000000000000000000, (if_mux_2_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_88_63 <= MUX_v_26_2_2(26'b00000000000000000000000000, (if_mux_3_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_114_89 <= MUX_v_26_2_2(26'b00000000000000000000000000, (if_mux_4_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_140_115 <= MUX_v_26_2_2(26'b00000000000000000000000000, (if_mux_5_nl),
          or_mdf_sva_mx0w0);
      hit_out_rsci_idat_141 <= (if_mux_6_nl) & or_mdf_sva_mx0w0;
      hit_out_rsci_idat_144_142 <= MUX_v_3_2_2(3'b000, (if_mux_7_nl), or_mdf_sva_mx0w0);
      hit_out_rsci_idat_171_145 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (if_mux_8_nl), or_mdf_sva_mx0w0);
      hit_out_rsci_idat_198_172 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (if_mux_9_nl), or_mdf_sva_mx0w0);
      hit_out_rsci_idat_225_199 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (if_mux_10_nl), or_mdf_sva_mx0w0);
      reg_isHit_rsci_idat_cse <= or_mdf_sva_mx0w0;
      attenuation_chan_out_rsci_idat <= attenuation_chan_in_rsci_idat_mxwt;
      accumalated_color_chan_in_crt_sva <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_idat_26_0 <= 27'b000000000000000000000000000;
      accumalated_color_out_rsci_idat_53_27 <= 27'b000000000000000000000000000;
      accumalated_color_out_rsci_idat_80_54 <= 27'b000000000000000000000000000;
    end
    else if ( accumalated_color_out_and_cse ) begin
      accumalated_color_out_rsci_idat_26_0 <= mux_11_itm;
      accumalated_color_out_rsci_idat_53_27 <= mux_12_itm;
      accumalated_color_out_rsci_idat_80_54 <= MUX_v_27_2_2((accumalated_color_chan_in_crt_sva[80:54]),
          z_out, and_45_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_isHit_rsci_ivld_hit_psct_cse <= 1'b0;
      reg_accumalated_color_out_rsci_ivld_hit_psct_cse <= 1'b0;
      reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse <= 1'b0;
      else_mul_cmp_b <= 27'b000000000000000000000000000;
      else_mul_cmp_a <= 27'b000000000000000000000000000;
      params_in_crt_sva_64_38 <= 27'b000000000000000000000000000;
      attenuation_chan_in_crt_sva_53_27 <= 27'b000000000000000000000000000;
      mux_12_itm <= 27'b000000000000000000000000000;
    end
    else if ( hit_wen ) begin
      reg_isHit_rsci_ivld_hit_psct_cse <= fsm_output[1];
      reg_accumalated_color_out_rsci_ivld_hit_psct_cse <= fsm_output[5];
      reg_closest_so_far_outtwo_rsci_irdy_hit_psct_cse <= (fsm_output[0]) | (fsm_output[6]);
      else_mul_cmp_b <= MUX1HOT_v_27_3_2((params_in_rsci_idat_mxwt[26:0]), params_in_crt_sva_64_38,
          params_in_crt_sva_91_65, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      else_mul_cmp_a <= MUX1HOT_v_27_3_2((attenuation_chan_in_rsci_idat_mxwt[26:0]),
          attenuation_chan_in_crt_sva_53_27, attenuation_chan_in_crt_sva_80_54, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[3])});
      params_in_crt_sva_64_38 <= params_in_rsci_idat_mxwt[53:27];
      attenuation_chan_in_crt_sva_53_27 <= attenuation_chan_in_rsci_idat_mxwt[53:27];
      mux_12_itm <= MUX_v_27_2_2(z_out, (accumalated_color_chan_in_crt_sva[53:27]),
          reg_isHit_rsci_idat_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_slc_47_svs <= 1'b0;
    end
    else if ( hit_wen & (~((~ (fsm_output[1])) | and_dcpl)) ) begin
      if_slc_47_svs <= if_acc_itm_47;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      params_in_crt_sva_91_65 <= 27'b000000000000000000000000000;
      attenuation_chan_in_crt_sva_80_54 <= 27'b000000000000000000000000000;
    end
    else if ( and_94_cse ) begin
      params_in_crt_sva_91_65 <= params_in_rsci_idat_mxwt[80:54];
      attenuation_chan_in_crt_sva_80_54 <= attenuation_chan_in_rsci_idat_mxwt[80:54];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mux_11_itm <= 27'b000000000000000000000000000;
    end
    else if ( hit_wen & (fsm_output[3]) ) begin
      mux_11_itm <= MUX_v_27_2_2((accumalated_color_chan_in_crt_sva[26:0]), z_out,
          and_82_nl);
    end
  end
  assign if_mux_nl = MUX_v_21_2_2((rec_quad_outtwo_rsci_idat_mxwt[20:0]), (rec_quad_outone_rsci_idat_mxwt[20:0]),
      if_acc_itm_47);
  assign if_mux_1_nl = MUX_v_21_2_2((rec_quad_outtwo_rsci_idat_mxwt[41:21]), (rec_quad_outone_rsci_idat_mxwt[41:21]),
      if_acc_itm_47);
  assign if_mux_2_nl = MUX_v_21_2_2((rec_quad_outtwo_rsci_idat_mxwt[62:42]), (rec_quad_outone_rsci_idat_mxwt[62:42]),
      if_acc_itm_47);
  assign if_mux_3_nl = MUX_v_26_2_2((rec_quad_outtwo_rsci_idat_mxwt[88:63]), (rec_quad_outone_rsci_idat_mxwt[88:63]),
      if_acc_itm_47);
  assign if_mux_4_nl = MUX_v_26_2_2((rec_quad_outtwo_rsci_idat_mxwt[114:89]), (rec_quad_outone_rsci_idat_mxwt[114:89]),
      if_acc_itm_47);
  assign if_mux_5_nl = MUX_v_26_2_2((rec_quad_outtwo_rsci_idat_mxwt[140:115]), (rec_quad_outone_rsci_idat_mxwt[140:115]),
      if_acc_itm_47);
  assign if_if_mux_1_nl = MUX_s_1_2_2(if_acc_itm_47, if_slc_47_svs, and_dcpl);
  assign if_mux_6_nl = MUX_s_1_2_2((rec_quad_outtwo_rsci_idat_mxwt[141]), (rec_quad_outone_rsci_idat_mxwt[141]),
      if_if_mux_1_nl);
  assign if_mux_7_nl = MUX_v_3_2_2((rec_quad_outtwo_rsci_idat_mxwt[144:142]), (rec_quad_outone_rsci_idat_mxwt[144:142]),
      if_acc_itm_47);
  assign if_mux_8_nl = MUX_v_27_2_2((rec_quad_outtwo_rsci_idat_mxwt[171:145]), (rec_quad_outone_rsci_idat_mxwt[171:145]),
      if_acc_itm_47);
  assign if_mux_9_nl = MUX_v_27_2_2((rec_quad_outtwo_rsci_idat_mxwt[198:172]), (rec_quad_outone_rsci_idat_mxwt[198:172]),
      if_acc_itm_47);
  assign if_mux_10_nl = MUX_v_27_2_2((rec_quad_outtwo_rsci_idat_mxwt[225:199]), (rec_quad_outone_rsci_idat_mxwt[225:199]),
      if_acc_itm_47);
  assign and_45_nl = (~ reg_isHit_rsci_idat_cse) & (fsm_output[5]);
  assign and_82_nl = (~ reg_isHit_rsci_idat_cse) & (fsm_output[3]);
  assign else_mux1h_3_nl = MUX1HOT_v_27_3_2((accumalated_color_chan_in_crt_sva[80:54]),
      (accumalated_color_chan_in_crt_sva[26:0]), (accumalated_color_chan_in_crt_sva[53:27]),
      {(fsm_output[5]) , (fsm_output[3]) , (fsm_output[4])});
  assign nl_z_out = else_mul_cmp_z_oreg + (else_mux1h_3_nl);
  assign z_out = nl_z_out[26:0];

  function automatic [26:0] MUX1HOT_v_27_3_2;
    input [26:0] input_2;
    input [26:0] input_1;
    input [26:0] input_0;
    input [2:0] sel;
    reg [26:0] result;
  begin
    result = input_0 & {27{sel[0]}};
    result = result | ( input_1 & {27{sel[1]}});
    result = result | ( input_2 & {27{sel[2]}});
    MUX1HOT_v_27_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_2_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input [0:0] sel;
    reg [25:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_26_2_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_2_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input [0:0] sel;
    reg [26:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_27_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_48_1_47;
    input [47:0] vector;
    reg [47:0] tmp;
  begin
    tmp = vector >> 47;
    readslicef_48_1_47 = tmp[0:0];
  end
  endfunction


  function automatic [47:0] conv_s2u_47_48 ;
    input [46:0]  vector ;
  begin
    conv_s2u_47_48 = {vector[46], vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter_scatter
// ------------------------------------------------------------------


module MaterialScatter_scatter (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, hit_in_rsc_dat, hit_in_rsc_vld,
      hit_in_rsc_rdy, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld, accumalated_color_chan_in_rsc_rdy,
      isHit_rsc_dat, isHit_rsc_vld, isHit_rsc_rdy, attenuation_chan_out_rsc_dat,
      attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy, accumalated_color_out_rsc_dat,
      accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy, ray_out_rsc_dat,
      ray_out_rsc_vld, ray_out_rsc_rdy, lambertianScatter_rand_unit_run_xs_mul_cmp_a,
      lambertianScatter_rand_unit_run_xs_mul_cmp_b, lambertianScatter_rand_unit_run_xs_mul_cmp_en,
      lambertianScatter_rand_unit_run_xs_mul_cmp_z, else_if_mul_cmp_a, else_if_mul_cmp_b,
      else_if_mul_cmp_z
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [225:0] hit_in_rsc_dat;
  input hit_in_rsc_vld;
  output hit_in_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input isHit_rsc_dat;
  input isHit_rsc_vld;
  output isHit_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  output [35:0] lambertianScatter_rand_unit_run_xs_mul_cmp_a;
  output [35:0] lambertianScatter_rand_unit_run_xs_mul_cmp_b;
  output lambertianScatter_rand_unit_run_xs_mul_cmp_en;
  input [65:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z;
  output [26:0] else_if_mul_cmp_a;
  reg [26:0] else_if_mul_cmp_a;
  output [26:0] else_if_mul_cmp_b;
  reg [26:0] else_if_mul_cmp_b;
  input [48:0] else_if_mul_cmp_z;


  // Interconnect Declarations
  wire scatter_wen;
  wire ray_in_rsci_wen_comp;
  wire [165:0] ray_in_rsci_idat_mxwt;
  wire hit_in_rsci_wen_comp;
  wire [225:0] hit_in_rsci_idat_mxwt;
  wire attenuation_chan_in_rsci_wen_comp;
  wire [80:0] attenuation_chan_in_rsci_idat_mxwt;
  wire accumalated_color_chan_in_rsci_wen_comp;
  wire [80:0] accumalated_color_chan_in_rsci_idat_mxwt;
  wire isHit_rsci_wen_comp;
  wire isHit_rsci_idat_mxwt;
  wire attenuation_chan_out_rsci_wen_comp;
  wire accumalated_color_out_rsci_wen_comp;
  wire ray_out_rsci_wen_comp;
  reg ensig_cgo;
  wire [33:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg;
  wire [26:0] else_if_mul_cmp_z_oreg;
  reg [26:0] attenuation_chan_out_rsci_idat_53_27;
  reg [26:0] accumalated_color_out_rsci_idat_80_54;
  reg [26:0] accumalated_color_out_rsci_idat_53_27;
  reg [26:0] accumalated_color_out_rsci_idat_26_0;
  reg ray_out_rsci_idat_165;
  reg [33:0] ray_out_rsci_idat_164_131;
  reg [33:0] ray_out_rsci_idat_130_97;
  reg [33:0] ray_out_rsci_idat_96_63;
  reg [20:0] ray_out_rsci_idat_62_42;
  reg [20:0] ray_out_rsci_idat_41_21;
  reg [20:0] ray_out_rsci_idat_20_0;
  wire [20:0] fsm_output;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_tmp;
  wire rand_unit_random2_run_x3_xor_26_tmp;
  wire and_dcpl_5;
  wire and_dcpl_18;
  wire or_dcpl_29;
  wire or_dcpl_30;
  wire or_dcpl_32;
  wire or_dcpl_35;
  wire or_dcpl_44;
  wire or_dcpl_45;
  wire and_dcpl_58;
  wire and_dcpl_62;
  wire or_dcpl_73;
  wire or_tmp_44;
  wire or_tmp_54;
  wire or_tmp_78;
  wire or_tmp_111;
  wire or_tmp_208;
  wire or_tmp_400;
  wire or_tmp_407;
  wire or_tmp_516;
  wire or_tmp_659;
  wire and_352_cse;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm;
  reg lambertianScatter_run_land_1_lpi_1_dfm;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_0;
  reg readHit_sva;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm;
  reg [63:0] ac_math_x2_acos_pi_2mi_64_return_sva;
  reg else_unequal_tmp;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1;
  reg rand_unit_random2_run_x3_31_sva;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42;
  reg [41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42;
  reg [41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0;
  reg [68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm;
  reg [1:0] reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd;
  reg [25:0] reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1;
  reg [7:0] reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2;
  reg [6:0] reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_3;
  reg [25:0] reg_lambertianScatter_add_run_acc_3_psp_ftd;
  reg [25:0] reg_lambertianScatter_add_run_acc_psp_ftd;
  wire ray_out_and_cse;
  wire accumalated_color_out_and_cse;
  reg reg_ray_out_rsci_ivld_scatter_psct_cse;
  reg reg_accumalated_color_out_rsci_ivld_scatter_psct_cse;
  reg reg_isHit_rsci_irdy_scatter_psct_cse;
  wire lambertianScatter_state1_and_cse;
  reg reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_1_2_svs_cse;
  reg reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_acc_1_2_svs_cse;
  wire else_and_cse;
  wire nor_cse;
  wire and_8_cse;
  reg rand_unit_random1_run_x3_sva_31;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva;
  wire ensig_cgo_mx0;
  reg rand_unit_random1_run_x3_sva_30;
  reg rand_unit_random1_run_x3_sva_29;
  reg rand_unit_random1_run_x3_sva_28;
  reg rand_unit_random1_run_x3_sva_27;
  reg rand_unit_random1_run_x3_sva_26;
  reg rand_unit_random1_run_x3_sva_25;
  reg rand_unit_random1_run_x3_sva_24;
  reg rand_unit_random1_run_x3_sva_23;
  reg rand_unit_random1_run_x3_sva_22;
  reg rand_unit_random1_run_x3_sva_21;
  reg rand_unit_random1_run_x3_sva_20;
  reg rand_unit_random1_run_x3_sva_19;
  reg rand_unit_random1_run_x3_sva_18;
  reg rand_unit_random1_run_x3_sva_17;
  reg rand_unit_random1_run_x3_sva_16;
  reg rand_unit_random1_run_x3_sva_15;
  reg rand_unit_random1_run_x3_sva_14;
  reg rand_unit_random1_run_x3_sva_13;
  reg rand_unit_random1_run_x3_sva_12;
  reg rand_unit_random1_run_x3_sva_11;
  reg rand_unit_random1_run_x3_sva_10;
  reg rand_unit_random1_run_x3_sva_9;
  reg rand_unit_random1_run_x3_sva_8;
  reg rand_unit_random1_run_x3_sva_7;
  reg rand_unit_random1_run_x3_sva_6;
  reg rand_unit_random1_run_x3_sva_5;
  reg rand_unit_random1_run_x2_12_0_sva_4;
  reg rand_unit_random1_run_x2_12_0_sva_3;
  reg rand_unit_random1_run_x2_12_0_sva_2;
  reg rand_unit_random1_run_x2_12_0_sva_1;
  reg rand_unit_random1_run_x2_12_0_sva_0;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_else_if_mux_1_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_mux_1_cse;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_itm;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_itm;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_itm;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_itm;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_itm;
  wire [42:0] operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm;
  wire [26:0] z_out;
  wire [27:0] nl_z_out;
  wire [31:0] z_out_3;
  wire [32:0] nl_z_out_3;
  wire [28:0] z_out_4;
  wire [29:0] nl_z_out_4;
  wire or_tmp_1118;
  wire or_tmp_1119;
  wire [69:0] z_out_5;
  wire [45:0] z_out_6;
  wire [45:0] z_out_7;
  wire [45:0] z_out_8;
  wire [45:0] z_out_9;
  wire [42:0] z_out_10;
  wire [42:0] z_out_11;
  wire [42:0] z_out_12;
  wire [42:0] z_out_13;
  wire [42:0] z_out_14;
  wire [42:0] z_out_15;
  wire [42:0] z_out_16;
  wire [42:0] z_out_17;
  wire [26:0] z_out_18;
  wire [27:0] nl_z_out_18;
  wire [68:0] z_out_19;
  wire [68:0] z_out_20;
  reg lambertianScatter_state2_15_sva;
  reg lambertianScatter_state2_16_sva;
  reg lambertianScatter_state2_14_sva;
  reg lambertianScatter_state2_17_sva;
  reg lambertianScatter_state2_13_sva;
  reg lambertianScatter_state2_18_sva;
  reg lambertianScatter_state2_12_sva;
  reg lambertianScatter_state2_19_sva;
  reg lambertianScatter_state2_11_sva;
  reg lambertianScatter_state2_20_sva;
  reg lambertianScatter_state2_10_sva;
  reg lambertianScatter_state2_21_sva;
  reg lambertianScatter_state2_9_sva;
  reg lambertianScatter_state2_22_sva;
  reg lambertianScatter_state2_8_sva;
  reg lambertianScatter_state2_23_sva;
  reg lambertianScatter_state2_7_sva;
  reg lambertianScatter_state2_24_sva;
  reg lambertianScatter_state2_6_sva;
  reg lambertianScatter_state2_25_sva;
  reg lambertianScatter_state2_5_sva;
  reg lambertianScatter_state2_26_sva;
  reg lambertianScatter_state2_4_sva;
  reg lambertianScatter_state2_27_sva;
  reg lambertianScatter_state2_3_sva;
  reg lambertianScatter_state2_28_sva;
  reg lambertianScatter_state2_2_sva;
  reg lambertianScatter_state2_29_sva;
  reg lambertianScatter_state2_1_sva;
  reg lambertianScatter_state2_30_sva;
  reg lambertianScatter_state2_0_sva;
  reg lambertianScatter_state2_31_sva;
  reg [165:0] ray_in_crt_sva;
  reg [80:0] accumalated_color_chan_in_crt_sva;
  reg [68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva;
  reg [68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva;
  reg [68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_sva;
  reg [68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva;
  wire [70:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva;
  reg [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva;
  reg [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva;
  reg [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva;
  reg [41:0] ac_math_atan_pi_2mi_return_69_28_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_2mi_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_sva;
  reg [41:0] ac_math_atan_pi_2mi_return_1_69_28_sva;
  reg [41:0] ac_math_atan_pi_2mi_return_2_69_28_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_x_2mi_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_y_2mi_sva;
  reg [41:0] ac_math_atan_pi_2mi_return_3_69_28_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_x_2mi_sva;
  reg [42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_y_2mi_sva;
  reg [26:0] lambertianScatter_add_run_acc_4_psp_sva;
  reg [20:0] mux_21_itm;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_42_39;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_38;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_37_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_29_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_25;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_24_23;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_22_20;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_10;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_9_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_5;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_4_1;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_0;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_42_39;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_38;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_35_34;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_33;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_32_31;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_30;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_29_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_25;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_22_20;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_18_17;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_16;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_15_14;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_10;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_5;
  reg [4:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_4_0;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_38;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_9_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_5;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_42_39;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_35_34;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_32_31;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_29_27;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_22_20;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14;
  reg [4:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_4_0;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_42_39;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_38;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_37_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_25;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_24_23;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_10;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_9_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_5;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_4_1;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_0;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_42_39;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_35_34;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_32_31;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_29_27;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_22_20;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_18_17;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_15_14;
  reg [4:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_4_0;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_42_39;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_38;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_37_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_29_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_25;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_24_23;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_10;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_9_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_5;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_4_1;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_0;
  reg [3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_42_39;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_38;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_35_34;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_33;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_32_31;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_30;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_29_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_25;
  reg [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_22_20;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_19;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_18_17;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_16;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_15_14;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_10;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_5;
  reg [4:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_4_0;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_35_34;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_32_31;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_18_17;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_35_34;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_32_31;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_15_14;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_38;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_33;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_30;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_26;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_25;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_19;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_16;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_13;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_12;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_11;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_10;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_5;
  reg lambertianScatter_state1_sva_31;
  reg lambertianScatter_state1_sva_30;
  reg lambertianScatter_state1_sva_29;
  reg lambertianScatter_state1_sva_28;
  reg lambertianScatter_state1_sva_27;
  reg lambertianScatter_state1_sva_26;
  reg lambertianScatter_state1_sva_25;
  reg lambertianScatter_state1_sva_24;
  reg lambertianScatter_state1_sva_23;
  reg lambertianScatter_state1_sva_22;
  reg lambertianScatter_state1_sva_21;
  reg lambertianScatter_state1_sva_20;
  reg lambertianScatter_state1_sva_19;
  reg lambertianScatter_state1_sva_18;
  reg lambertianScatter_state1_sva_17;
  reg lambertianScatter_state1_sva_16;
  reg lambertianScatter_state1_sva_15;
  reg lambertianScatter_state1_sva_14;
  reg lambertianScatter_state1_sva_13;
  reg lambertianScatter_state1_sva_12;
  reg lambertianScatter_state1_sva_11;
  reg lambertianScatter_state1_sva_10;
  reg lambertianScatter_state1_sva_9;
  reg lambertianScatter_state1_sva_8;
  reg lambertianScatter_state1_sva_7;
  reg lambertianScatter_state1_sva_6;
  reg lambertianScatter_state1_sva_5;
  reg lambertianScatter_state1_sva_4;
  reg lambertianScatter_state1_sva_3;
  reg lambertianScatter_state1_sva_2;
  reg lambertianScatter_state1_sva_1;
  reg lambertianScatter_state1_sva_0;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0;
  reg [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_37;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_24;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_23;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_9;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_8;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_7;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_29;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_29;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_28;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_27;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_22;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_21;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_20;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_37;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_24;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_23;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_9;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_8;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_7;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_37;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_36;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_24;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_23;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_9;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_8;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_7;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_6;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_35;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_34;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_32;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_31;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_18;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_17;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_15;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_14;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_35;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_34;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_32;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_31;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_18;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_17;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_15;
  reg ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_14;
  wire rand_unit_random2_run_x3_11_sva_mx0w0;
  wire rand_unit_random2_run_x2_1_sva_mx0w0;
  wire rand_unit_random2_run_x3_10_sva_mx0w0;
  wire rand_unit_random2_run_x2_0_sva_mx0w0;
  wire rand_unit_random2_run_x2_4_sva_mx0w0;
  wire rand_unit_random2_run_x2_3_sva_mx0w0;
  wire rand_unit_random2_run_x2_2_sva_mx0w0;
  wire rand_unit_random2_run_x3_17_sva_mx0w0;
  wire rand_unit_random2_run_x3_28_sva_mx0w0;
  wire rand_unit_random2_run_x3_9_sva_mx0w0;
  wire rand_unit_random2_run_x3_5_sva_mx0w0;
  wire rand_unit_random2_run_x3_8_sva_mx0w0;
  wire rand_unit_random2_run_x3_6_sva_mx0w0;
  wire rand_unit_random2_run_x3_7_sva_mx0w0;
  wire rand_unit_random2_run_x3_30_sva_mx0w0;
  wire rand_unit_random2_run_x3_15_sva_mx0w0;
  wire rand_unit_random2_run_x3_14_sva_mx0w0;
  wire rand_unit_random2_run_x3_27_sva_mx0w0;
  wire rand_unit_random2_run_x3_13_sva_mx0w0;
  wire rand_unit_random2_run_x3_12_sva_mx0w0;
  wire rand_unit_random2_run_x3_26_sva_mx0w0;
  wire rand_unit_random2_run_x3_25_sva_mx0w0;
  wire rand_unit_random2_run_x3_24_sva_mx0w0;
  wire rand_unit_random2_run_x3_23_sva_mx0w0;
  wire rand_unit_random2_run_x3_16_sva_mx0w0;
  wire rand_unit_random2_run_x3_22_sva_mx0w0;
  wire rand_unit_random2_run_x3_18_sva_mx0w0;
  wire rand_unit_random2_run_x3_21_sva_mx0w0;
  wire rand_unit_random2_run_x3_19_sva_mx0w0;
  wire rand_unit_random2_run_x3_20_sva_mx0w0;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2;
  wire lambertianScatter_run_land_lpi_1_dfm_mx1w0;
  wire lambertianScatter_run_land_1_lpi_1_dfm_mx2;
  wire [64:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_lpi_1_dfm_64_0_mx0;
  wire [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1;
  wire [1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1;
  wire [2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1;
  wire [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3;
  wire [6:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3;
  wire [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2;
  wire [6:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2;
  wire [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1;
  wire [6:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1;
  wire [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2;
  wire [6:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs_mx0c2;
  wire [44:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6;
  wire [45:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6;
  wire [44:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6;
  wire [45:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6;
  wire [44:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6;
  wire [45:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6;
  wire [44:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6;
  wire [45:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6;
  wire xor_cse;
  wire xor_cse_1;
  wire xor_cse_2;
  wire xor_cse_3;
  wire xor_cse_4;
  wire xor_cse_5;
  wire xor_cse_6;
  wire xor_cse_7;
  wire xor_cse_8;
  wire xor_cse_9;
  wire xor_cse_10;
  wire xor_cse_11;
  wire xor_cse_12;
  wire xor_cse_13;
  wire xor_cse_14;
  wire xor_cse_15;
  wire xor_cse_16;
  wire xor_cse_17;
  wire xor_cse_18;
  wire xor_cse_19;
  wire xor_cse_20;
  wire xor_cse_21;
  wire xor_cse_22;
  wire xor_cse_23;
  wire xor_cse_24;
  wire xor_cse_25;
  wire xor_cse_26;
  wire xor_cse_27;
  wire xor_cse_28;
  wire xor_cse_29;
  wire xor_cse_30;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_theta_d_and_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_d_a_and_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_and_cse;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_1_ssc;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_4_ssc;
  reg [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36;
  reg [35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0;
  reg [5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36;
  reg [35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0;
  wire lambertianScatter_state2_and_32_cse;
  wire ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_45_cse;
  wire rand_unit_random2_run_x3_and_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_9_cse;
  reg reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_6_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_84_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_11_cse;
  wire [26:0] color_out_g_mux1h_5_rgt;
  wire [27:0] lambertianScatter_run_aelse_1_mux1h_7_rgt;
  wire [26:0] color_out_r_mux1h_3_rgt;
  wire and_dcpl_110;
  wire [65:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_rgt;
  wire [6:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_rgt;
  wire [6:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_rgt;
  wire [7:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_rgt;
  wire [32:0] lambertianScatter_rand_unit_run_phi_mux1h_2_rgt;
  reg ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65;
  reg [26:0] hit_in_crt_sva_198_172;
  reg [171:0] hit_in_crt_sva_171_0;
  reg [11:0] lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21;
  reg [20:0] lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0;
  reg lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_27;
  reg [26:0] lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0;
  reg [3:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_7_4;
  reg [3:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0;
  reg [2:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_6_4;
  reg [3:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0;
  reg [5:0] color_out_r_sva_1_26_21;
  reg [20:0] color_out_r_sva_1_20_0;
  reg color_out_g_sva_1_26;
  reg [25:0] color_out_g_sva_1_25_0;
  reg [26:0] attenuation_chan_in_crt_sva_53_27;
  reg [26:0] attenuation_chan_in_crt_sva_26_0;
  reg attenuation_chan_out_rsci_idat_80;
  reg [25:0] attenuation_chan_out_rsci_idat_79_54;
  reg [5:0] attenuation_chan_out_rsci_idat_26_21;
  reg [20:0] attenuation_chan_out_rsci_idat_20_0;
  wire or_1202_ssc;
  reg reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg;
  reg [5:0] reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg;
  reg [32:0] reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg;
  reg [31:0] reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg;
  wire color_out_g_and_1_cse;
  wire color_out_g_and_cse;
  wire and_2513_cse;
  wire and_2517_cse;
  wire and_2523_cse;
  wire and_2527_cse;
  wire nor_31_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_29_cse;
  wire and_2512_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_cse;
  wire ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_1_cse;
  wire z_out_1_33;
  wire z_out_21_2;

  wire[25:0] lambertianScatter_run_mux_nl;
  wire[25:0] lambertianScatter_run_mux_1_nl;
  wire[25:0] lambertianScatter_run_mux_2_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_4_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_8_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_17_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_41_nl;
  wire[6:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl;
  wire[7:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl;
  wire[26:0] color_out_b_color_out_b_mux_1_nl;
  wire[33:0] ac_math_ac_abs_35_35_xabs_acc_nl;
  wire[34:0] nl_ac_math_ac_abs_35_35_xabs_acc_nl;
  wire[33:0] ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_2_nl;
  wire[33:0] ac_math_ac_abs_35_35_xabs_xor_1_nl;
  wire[33:0] ac_math_ac_abs_35_35_2_xabs_xor_1_nl;
  wire[0:0] ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_3_nl;
  wire[0:0] and_945_nl;
  wire[0:0] lambertianScatter_run_aelse_1_or_nl;
  wire[20:0] hit_in_hit_loc_x_hit_in_hit_loc_x_mux_nl;
  wire[0:0] color_out_r_and_nl;
  wire[0:0] color_out_r_and_1_nl;
  wire[65:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_mux1h_4_nl;
  wire[65:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl;
  wire[67:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl;
  wire[65:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl;
  wire[66:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl;
  wire[0:0] not_343_nl;
  wire[6:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_nl;
  wire[5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_nl;
  wire[0:0] not_271_nl;
  wire[0:0] not_342_nl;
  wire[68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl;
  wire[70:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl;
  wire[68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl;
  wire[69:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl;
  wire[0:0] not_341_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_or_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_nor_nl;
  wire[3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_and_nl;
  wire[0:0] not_270_nl;
  wire[3:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_nl;
  wire[0:0] not_269_nl;
  wire[1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_5_nl;
  wire[0:0] not_340_nl;
  wire[1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_4_nl;
  wire[0:0] not_339_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux1h_89_nl;
  wire[32:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl;
  wire[33:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl;
  wire[20:0] hit_in_hit_loc_y_hit_in_hit_loc_y_mux_nl;
  wire[0:0] lambertianScatter_rand_unit_run_phi_and_nl;
  wire[0:0] lambertianScatter_rand_unit_run_phi_and_1_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_33_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_32_nl;
  wire[0:0] not_335_nl;
  wire[0:0] not_334_nl;
  wire[0:0] not_333_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_7_nl;
  wire[0:0] not_329_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_2_nl;
  wire[0:0] not_324_nl;
  wire[0:0] not_323_nl;
  wire[0:0] not_322_nl;
  wire[41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_1_nl;
  wire[0:0] not_321_nl;
  wire[0:0] not_320_nl;
  wire[5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_1_nl;
  wire[0:0] not_533_nl;
  wire[35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_16_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_or_3_nl;
  wire[0:0] and_202_nl;
  wire[0:0] not_319_nl;
  wire[0:0] not_318_nl;
  wire[0:0] not_317_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_6_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_5_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_4_nl;
  wire[0:0] not_313_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_3_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_2_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_1_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_nl;
  wire[0:0] not_308_nl;
  wire[0:0] not_307_nl;
  wire[5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_nl;
  wire[0:0] not_534_nl;
  wire[35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_15_nl;
  wire[0:0] and_204_nl;
  wire[0:0] not_306_nl;
  wire[0:0] not_305_nl;
  wire[41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_nl;
  wire[0:0] not_304_nl;
  wire[0:0] not_303_nl;
  wire[0:0] not_302_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_10_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl;
  wire[0:0] not_298_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_6_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl;
  wire[0:0] not_293_nl;
  wire[0:0] not_292_nl;
  wire[0:0] else_else_and_1_nl;
  wire[0:0] lambertianScatter_run_if_lambertianScatter_run_if_and_1_nl;
  wire[64:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[65:0] nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[6:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl;
  wire[7:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl;
  wire[6:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl;
  wire[7:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl;
  wire[6:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl;
  wire[7:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl;
  wire[6:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl;
  wire[7:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl;
  wire[26:0] else_else_mux1h_1_nl;
  wire[33:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl;
  wire[34:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_32_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_33_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_34_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_35_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_36_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_37_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_38_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_39_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_40_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_41_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_42_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_43_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_44_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_45_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_46_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_47_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_48_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_49_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_50_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_51_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_52_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_53_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_54_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_55_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_56_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_57_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_58_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_59_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_60_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_61_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_62_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_63_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_nand_1_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_31_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_31_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_32_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_33_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_32_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_34_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_33_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_35_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_34_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_36_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_35_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_37_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_36_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_38_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_37_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_39_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_38_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_40_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_39_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_41_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_40_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_42_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_41_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_43_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_42_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_44_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_43_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_45_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_44_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_46_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_45_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_47_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_46_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_48_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_47_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_49_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_48_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_50_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_49_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_51_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_50_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_52_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_51_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_53_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_52_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_54_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_53_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_55_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_54_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_56_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_55_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_57_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_56_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_58_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_57_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_59_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_58_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_60_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_59_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_61_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_60_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_2_nl;
  wire[19:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_3_nl;
  wire[6:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_2_nl;
  wire[70:0] acc_5_nl;
  wire[71:0] nl_acc_5_nl;
  wire[68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_1_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_4_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_5_nl;
  wire[68:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux1h_1_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_6_nl;
  wire[0:0] ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_7_nl;
  wire[46:0] acc_6_nl;
  wire[47:0] nl_acc_6_nl;
  wire[2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_33_nl;
  wire[5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_34_nl;
  wire[35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_35_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_36_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_37_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_38_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_39_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_40_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_41_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_42_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_43_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_44_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_45_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_46_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_47_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_48_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_49_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_50_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_51_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_52_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_53_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_54_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_55_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_56_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_57_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_58_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_59_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_60_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_61_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_62_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_63_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_64_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_65_nl;
  wire[11:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_n000000;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_not_61_nl;
  wire[46:0] acc_7_nl;
  wire[47:0] nl_acc_7_nl;
  wire[2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_32_nl;
  wire[41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_33_nl;
  wire[43:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_34_nl;
  wire[46:0] acc_8_nl;
  wire[47:0] nl_acc_8_nl;
  wire[2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_63_nl;
  wire[5:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_64_nl;
  wire[35:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_65_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_66_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_67_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_68_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_69_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_70_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_71_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_72_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_73_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_74_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_75_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_76_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_77_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_78_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_79_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_80_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_81_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_82_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_83_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_84_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_85_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_86_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_87_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_88_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_89_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_90_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_91_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_92_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_93_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_94_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_95_nl;
  wire[11:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_n000000;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_not_61_nl;
  wire[46:0] acc_9_nl;
  wire[47:0] nl_acc_9_nl;
  wire[2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_32_nl;
  wire[41:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_33_nl;
  wire[43:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_34_nl;
  wire[43:0] acc_10_nl;
  wire[44:0] nl_acc_10_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_nand_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_mux_29_nl;
  wire[43:0] acc_11_nl;
  wire[44:0] nl_acc_11_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_nand_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_35_nl;
  wire[43:0] acc_12_nl;
  wire[44:0] nl_acc_12_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_29_nl;
  wire[43:0] acc_13_nl;
  wire[44:0] nl_acc_13_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_or_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_96_nl;
  wire[43:0] acc_14_nl;
  wire[44:0] nl_acc_14_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_nand_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_mux_29_nl;
  wire[43:0] acc_15_nl;
  wire[44:0] nl_acc_15_nl;
  wire[3:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_29_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_30_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_31_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_32_nl;
  wire[1:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_33_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_34_nl;
  wire[1:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_35_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_36_nl;
  wire[2:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_37_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_38_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_39_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_40_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_41_nl;
  wire[2:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_42_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_43_nl;
  wire[1:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_44_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_45_nl;
  wire[1:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_46_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_47_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_48_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_49_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_50_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_51_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_52_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_53_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_54_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_55_nl;
  wire[4:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_56_nl;
  wire[0:0] lambertianScatter_add_run_or_30_nl;
  wire[1:0] lambertianScatter_add_run_mux1h_44_nl;
  wire[0:0] lambertianScatter_add_run_lambertianScatter_add_run_mux_57_nl;
  wire[24:0] lambertianScatter_add_run_mux1h_45_nl;
  wire[7:0] lambertianScatter_add_run_mux1h_46_nl;
  wire[6:0] lambertianScatter_add_run_mux1h_47_nl;
  wire[43:0] acc_16_nl;
  wire[44:0] nl_acc_16_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_or_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_mux_29_nl;
  wire[43:0] acc_17_nl;
  wire[44:0] nl_acc_17_nl;
  wire[0:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_or_1_nl;
  wire[42:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_35_nl;
  wire[25:0] lambertianScatter_add_run_mux_8_nl;
  wire[2:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl;
  wire[3:0] nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl;
  wire[1:0] ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_a = {ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_29
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_22
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_21
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_0};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_s = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva;
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_a = {ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_4_0};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_s = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva;
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_4_0};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_s = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva;
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_a = {ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_4_0};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_s = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva;
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_a = {ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_35
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_32
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_18
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_15
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_0};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_s = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva;
  wire [42:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_a = {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_29
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_18_17
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_5
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12};
  wire [5:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_s = reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg;
  wire [68:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_a = MUX1HOT_v_69_3_2(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva,
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm,
      (signext_69_43({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_4_0})),
      {(fsm_output[6]) , (fsm_output[7]) , (fsm_output[12])});
  wire [7:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_s;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_s = MUX1HOT_v_8_3_2((z_out_4[7:0]),
      ({ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_7_4
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0}),
      ({2'b00 , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg}),
      {(fsm_output[6]) , (fsm_output[7]) , (fsm_output[12])});
  wire [68:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_a = MUX1HOT_v_69_4_2((~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva),
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva, (~
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm),
      (signext_69_43({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_35
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_32
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_18
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_15
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_0})),
      {(fsm_output[7]) , (fsm_output[8]) , (fsm_output[6]) , (fsm_output[12])});
  wire[0:0] operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl;
  wire[0:0] operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_1_nl;
  wire[4:0] operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_mux_nl;
  wire[0:0] operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl;
  wire [7:0] nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl
      = reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg
      & (~ (fsm_output[12]));
  assign operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_1_nl
      = (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[5])
      & (~ (fsm_output[12]));
  assign operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_mux_nl
      = MUX_v_5_2_2((reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[4:0]),
      (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva[5:1]),
      fsm_output[12]);
  assign operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl
      = (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva[0])
      & (fsm_output[8:6]==3'b000);
  assign nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_s = {(operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl)
      , (operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_1_nl)
      , (operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_mux_nl)
      , (operator_69_3_true_AC_TRN_AC_WRAP_3_operator_69_3_true_AC_TRN_AC_WRAP_3_and_nl)};
  wire [80:0] nl_MaterialScatter_scatter_attenuation_chan_out_rsci_inst_attenuation_chan_out_rsci_idat;
  assign nl_MaterialScatter_scatter_attenuation_chan_out_rsci_inst_attenuation_chan_out_rsci_idat
      = {attenuation_chan_out_rsci_idat_80 , attenuation_chan_out_rsci_idat_79_54
      , attenuation_chan_out_rsci_idat_53_27 , attenuation_chan_out_rsci_idat_26_21
      , attenuation_chan_out_rsci_idat_20_0};
  wire [80:0] nl_MaterialScatter_scatter_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat;
  assign nl_MaterialScatter_scatter_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat
      = {accumalated_color_out_rsci_idat_80_54 , accumalated_color_out_rsci_idat_53_27
      , accumalated_color_out_rsci_idat_26_0};
  wire [165:0] nl_MaterialScatter_scatter_ray_out_rsci_inst_ray_out_rsci_idat;
  assign nl_MaterialScatter_scatter_ray_out_rsci_inst_ray_out_rsci_idat = {ray_out_rsci_idat_165
      , ray_out_rsci_idat_164_131 , ray_out_rsci_idat_130_97 , ray_out_rsci_idat_96_63
      , ray_out_rsci_idat_62_42 , ray_out_rsci_idat_41_21 , ray_out_rsci_idat_20_0};
  wire [0:0] nl_MaterialScatter_scatter_scatter_fsm_inst_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0;
  assign nl_MaterialScatter_scatter_scatter_fsm_inst_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0
      = ~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm;
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd43),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd43)) operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_a[42:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_rg_s[5:0]),
      .z(operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd69),
  .signd_a(32'sd1),
  .width_s(32'sd8),
  .width_z(32'sd69)) operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_a[68:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_3_rshift_rg_s[7:0]),
      .z(z_out_19)
    );
  mgc_shift_r_v5 #(.width_a(32'sd69),
  .signd_a(32'sd1),
  .width_s(32'sd8),
  .width_z(32'sd69)) operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_a[68:0]),
      .s(nl_operator_43_4_true_AC_TRN_AC_WRAP_rshift_rg_s[7:0]),
      .z(z_out_20)
    );
  MaterialScatter_scatter_ray_in_rsci MaterialScatter_scatter_ray_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .scatter_wen(scatter_wen),
      .ray_in_rsci_oswt(reg_isHit_rsci_irdy_scatter_psct_cse),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .ray_in_rsci_idat_mxwt(ray_in_rsci_idat_mxwt)
    );
  MaterialScatter_scatter_hit_in_rsci MaterialScatter_scatter_hit_in_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .hit_in_rsc_dat(hit_in_rsc_dat),
      .hit_in_rsc_vld(hit_in_rsc_vld),
      .hit_in_rsc_rdy(hit_in_rsc_rdy),
      .scatter_wen(scatter_wen),
      .hit_in_rsci_oswt(reg_isHit_rsci_irdy_scatter_psct_cse),
      .hit_in_rsci_wen_comp(hit_in_rsci_wen_comp),
      .hit_in_rsci_idat_mxwt(hit_in_rsci_idat_mxwt)
    );
  MaterialScatter_scatter_attenuation_chan_in_rsci MaterialScatter_scatter_attenuation_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .scatter_wen(scatter_wen),
      .attenuation_chan_in_rsci_oswt(reg_isHit_rsci_irdy_scatter_psct_cse),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_idat_mxwt(attenuation_chan_in_rsci_idat_mxwt)
    );
  MaterialScatter_scatter_accumalated_color_chan_in_rsci MaterialScatter_scatter_accumalated_color_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .scatter_wen(scatter_wen),
      .accumalated_color_chan_in_rsci_oswt(reg_isHit_rsci_irdy_scatter_psct_cse),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_idat_mxwt(accumalated_color_chan_in_rsci_idat_mxwt)
    );
  MaterialScatter_scatter_isHit_rsci MaterialScatter_scatter_isHit_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .isHit_rsc_dat(isHit_rsc_dat),
      .isHit_rsc_vld(isHit_rsc_vld),
      .isHit_rsc_rdy(isHit_rsc_rdy),
      .scatter_wen(scatter_wen),
      .isHit_rsci_oswt(reg_isHit_rsci_irdy_scatter_psct_cse),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp),
      .isHit_rsci_idat_mxwt(isHit_rsci_idat_mxwt)
    );
  MaterialScatter_scatter_attenuation_chan_out_rsci MaterialScatter_scatter_attenuation_chan_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .scatter_wen(scatter_wen),
      .attenuation_chan_out_rsci_oswt(reg_accumalated_color_out_rsci_ivld_scatter_psct_cse),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .attenuation_chan_out_rsci_idat(nl_MaterialScatter_scatter_attenuation_chan_out_rsci_inst_attenuation_chan_out_rsci_idat[80:0])
    );
  MaterialScatter_scatter_accumalated_color_out_rsci MaterialScatter_scatter_accumalated_color_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .scatter_wen(scatter_wen),
      .accumalated_color_out_rsci_oswt(reg_accumalated_color_out_rsci_ivld_scatter_psct_cse),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .accumalated_color_out_rsci_idat(nl_MaterialScatter_scatter_accumalated_color_out_rsci_inst_accumalated_color_out_rsci_idat[80:0])
    );
  MaterialScatter_scatter_ray_out_rsci MaterialScatter_scatter_ray_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .scatter_wen(scatter_wen),
      .ray_out_rsci_oswt(reg_ray_out_rsci_ivld_scatter_psct_cse),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_idat(nl_MaterialScatter_scatter_ray_out_rsci_inst_ray_out_rsci_idat[165:0])
    );
  MaterialScatter_scatter_wait_dp MaterialScatter_scatter_wait_dp_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ensig_cgo_iro(ensig_cgo_mx0),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_en(lambertianScatter_rand_unit_run_xs_mul_cmp_en),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_z(lambertianScatter_rand_unit_run_xs_mul_cmp_z),
      .else_if_mul_cmp_z(else_if_mul_cmp_z),
      .scatter_wen(scatter_wen),
      .ensig_cgo(ensig_cgo),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg(lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg),
      .else_if_mul_cmp_z_oreg(else_if_mul_cmp_z_oreg)
    );
  MaterialScatter_scatter_staller MaterialScatter_scatter_staller_inst (
      .scatter_wen(scatter_wen),
      .ray_in_rsci_wen_comp(ray_in_rsci_wen_comp),
      .hit_in_rsci_wen_comp(hit_in_rsci_wen_comp),
      .attenuation_chan_in_rsci_wen_comp(attenuation_chan_in_rsci_wen_comp),
      .accumalated_color_chan_in_rsci_wen_comp(accumalated_color_chan_in_rsci_wen_comp),
      .isHit_rsci_wen_comp(isHit_rsci_wen_comp),
      .attenuation_chan_out_rsci_wen_comp(attenuation_chan_out_rsci_wen_comp),
      .accumalated_color_out_rsci_wen_comp(accumalated_color_out_rsci_wen_comp),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp)
    );
  MaterialScatter_scatter_scatter_fsm MaterialScatter_scatter_scatter_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .scatter_wen(scatter_wen),
      .fsm_output(fsm_output),
      .main_C_4_tr0(or_dcpl_30),
      .ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0(nl_MaterialScatter_scatter_scatter_fsm_inst_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_2_tr0[0:0]),
      .main_C_7_tr0(or_dcpl_30),
      .ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_C_1_tr0(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm)
    );
  assign ray_out_and_cse = scatter_wen & (fsm_output[19]);
  assign accumalated_color_out_and_cse = scatter_wen & (fsm_output[14]);
  assign lambertianScatter_state2_and_32_cse = scatter_wen & (~ else_unequal_tmp)
      & or_tmp_78;
  assign lambertianScatter_state1_and_cse = scatter_wen & ((isHit_rsci_idat_mxwt
      & (hit_in_rsci_idat_mxwt[144:142]==3'b000) & (fsm_output[1])) | or_tmp_111);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
      = (~ rand_unit_random2_run_x3_xor_26_tmp) & (fsm_output[1]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
      = rand_unit_random2_run_x3_xor_26_tmp & (fsm_output[1]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_45_cse
      = scatter_wen & (~ or_tmp_208);
  assign rand_unit_random2_run_x3_and_cse = scatter_wen & (~(and_dcpl_62 & and_dcpl_58
      & (~ (fsm_output[16])) & (~ (fsm_output[14]))));
  assign else_and_cse = scatter_wen & (fsm_output[1]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse
      = (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1)
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_84_cse
      = scatter_wen & (~(or_dcpl_45 | (fsm_output[4]) | (fsm_output[11]) | (fsm_output[12])));
  assign color_out_g_and_1_cse = else_unequal_tmp & (fsm_output[4]);
  assign color_out_g_mux1h_5_rgt = MUX1HOT_v_27_3_2(else_if_mul_cmp_z_oreg, z_out,
      ({1'b0 , (hit_in_crt_sva_171_0[114:89])}), {(fsm_output[3]) , color_out_g_and_1_cse
      , or_dcpl_32});
  assign color_out_g_and_cse = (~ else_unequal_tmp) & (fsm_output[4]);
  assign color_out_b_color_out_b_mux_1_nl = MUX_v_27_2_2(z_out, else_if_mul_cmp_z_oreg,
      color_out_g_and_cse);
  assign ac_math_ac_abs_35_35_xabs_xor_1_nl = (signext_34_1(z_out_18[26])) ^ ({(z_out_18[25:0])
      , (lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg[7:0])});
  assign ac_math_ac_abs_35_35_2_xabs_xor_1_nl = (signext_34_1(lambertianScatter_add_run_acc_4_psp_sva[26]))
      ^ ({(lambertianScatter_add_run_acc_4_psp_sva[25:0]) , reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2});
  assign ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_2_nl = MUX_v_34_2_2((ac_math_ac_abs_35_35_xabs_xor_1_nl),
      (ac_math_ac_abs_35_35_2_xabs_xor_1_nl), fsm_output[18]);
  assign ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_3_nl = MUX_s_1_2_2((z_out_18[26]),
      (lambertianScatter_add_run_acc_4_psp_sva[26]), fsm_output[18]);
  assign nl_ac_math_ac_abs_35_35_xabs_acc_nl = (ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_2_nl)
      + conv_u2u_1_34(ac_math_ac_abs_35_35_xabs_ac_math_ac_abs_35_35_xabs_mux_3_nl);
  assign ac_math_ac_abs_35_35_xabs_acc_nl = nl_ac_math_ac_abs_35_35_xabs_acc_nl[33:0];
  assign and_945_nl = and_dcpl_62 & and_dcpl_58 & (~ (fsm_output[16])) & (~ (fsm_output[2]))
      & (~ (fsm_output[14]));
  assign lambertianScatter_run_aelse_1_or_nl = (fsm_output[18:16]!=3'b000);
  assign lambertianScatter_run_aelse_1_mux1h_7_rgt = MUX1HOT_v_28_3_2(({1'b0 , (color_out_b_color_out_b_mux_1_nl)}),
      ({2'b00 , (hit_in_crt_sva_171_0[88:63])}), (readslicef_34_28_6((ac_math_ac_abs_35_35_xabs_acc_nl))),
      {(and_945_nl) , (fsm_output[15]) , (lambertianScatter_run_aelse_1_or_nl)});
  assign nor_31_cse = ~((fsm_output[20]) | (fsm_output[0]));
  assign hit_in_hit_loc_x_hit_in_hit_loc_x_mux_nl = MUX_v_21_2_2((hit_in_crt_sva_171_0[20:0]),
      (ray_in_crt_sva[20:0]), and_352_cse);
  assign color_out_r_and_nl = (~ else_unequal_tmp) & (fsm_output[5]);
  assign color_out_r_and_1_nl = else_unequal_tmp & (fsm_output[5]);
  assign color_out_r_mux1h_3_rgt = MUX1HOT_v_27_3_2(else_if_mul_cmp_z_oreg, z_out,
      ({6'b000000 , (hit_in_hit_loc_x_hit_in_hit_loc_x_mux_nl)}), {(color_out_r_and_nl)
      , (color_out_r_and_1_nl) , or_tmp_400});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
      & (fsm_output[7]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse
      = (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1)
      & (fsm_output[7]);
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl
      = ({ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg})
      + conv_s2s_65_66({1'b1 , (~ ac_math_x2_acos_pi_2mi_64_return_sva)}) + 66'b000000000000000000000000000000000000000000000000000000000000000001;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl[65:0];
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl
      = ({ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg})
      + conv_u2s_64_66(ac_math_x2_acos_pi_2mi_64_return_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl[65:0];
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_mux1h_4_nl
      = MUX1HOT_v_66_3_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_acc_2_nl),
      (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_acc_2_nl),
      ({1'b0 , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_lpi_1_dfm_64_0_mx0[64:32])
      , 32'b00000000000000000000000000000000}), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse
      , (fsm_output[9])});
  assign not_343_nl = ~ (fsm_output[5]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_rgt
      = MUX_v_66_2_2(66'b000000000000000000000000000000000000000000000000000000000000000000,
      (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_mux1h_4_nl),
      (not_343_nl));
  assign not_271_nl = ~ or_tmp_659;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_nl
      = MUX_v_6_2_2(6'b000000, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1,
      (not_271_nl));
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_nl
      = MUX_v_7_2_2(({ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_6_4
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0}),
      ({1'b0 , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_nl)}),
      or_tmp_407);
  assign not_342_nl = ~ (fsm_output[5]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_rgt
      = MUX_v_7_2_2(7'b0000000, (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_nl),
      (not_342_nl));
  assign and_8_cse = (~ else_unequal_tmp) & readHit_sva;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_theta_d_and_cse
      = scatter_wen & nor_cse & (~ (hit_in_crt_sva_171_0[142])) & readHit_sva;
  assign not_270_nl = ~ or_tmp_659;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_and_nl
      = MUX_v_4_2_2(4'b0000, (z_out_14[42:39]), (not_270_nl));
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_rgt
      = MUX_v_7_2_2((z_out_3[6:0]), ({3'b000 , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_else_and_nl)}),
      or_tmp_407);
  assign not_269_nl = ~ or_tmp_659;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_nl
      = MUX_v_4_2_2(4'b0000, (z_out_14[4:1]), (not_269_nl));
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_rgt
      = MUX_v_8_2_2((z_out_4[7:0]), ({4'b0000 , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_nl)}),
      or_tmp_407);
  assign and_2512_cse = (~ (fsm_output[12])) & scatter_wen;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_9_cse
      = scatter_wen & (fsm_output[12:10]==3'b000);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_29_cse
      = scatter_wen & (~ (fsm_output[10]));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse
      = (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs)
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse;
  assign and_2513_cse = ((fsm_output[13]) | (fsm_output[9]) | (fsm_output[11])) &
      scatter_wen;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_6_cse
      = scatter_wen & (~ or_tmp_516);
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl
      = (~ reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg)
      + ({32'b10000000000000000000000000000000 , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl[32:0];
  assign hit_in_hit_loc_y_hit_in_hit_loc_y_mux_nl = MUX_v_21_2_2((hit_in_crt_sva_171_0[41:21]),
      (ray_in_crt_sva[41:21]), and_352_cse);
  assign lambertianScatter_rand_unit_run_phi_and_nl = (~ rand_unit_random2_run_x3_31_sva)
      & (fsm_output[10]);
  assign lambertianScatter_rand_unit_run_phi_and_1_nl = rand_unit_random2_run_x3_31_sva
      & (fsm_output[10]);
  assign lambertianScatter_rand_unit_run_phi_mux1h_2_rgt = MUX1HOT_v_33_3_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_acc_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg,
      ({12'b000000000000 , (hit_in_hit_loc_y_hit_in_hit_loc_y_mux_nl)}), {(lambertianScatter_rand_unit_run_phi_and_nl)
      , (lambertianScatter_rand_unit_run_phi_and_1_nl) , or_tmp_400});
  assign and_2517_cse = ((fsm_output[13]) | (fsm_output[11])) & scatter_wen;
  assign and_2523_cse = (~ (fsm_output[13])) & scatter_wen;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt
      = (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs)
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_4_ssc
      = (~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs))
      & (fsm_output[13]);
  assign and_2527_cse = (((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm)
      & (fsm_output[13])) | (fsm_output[11])) & scatter_wen;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_11_cse
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_1_ssc
      = (~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm
      | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1))
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt
      = (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs)
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_d_a_and_cse
      = scatter_wen & (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_tmp);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_and_cse
      = scatter_wen & and_dcpl_5 & and_dcpl_18;
  assign nor_cse = ~((hit_in_crt_sva_171_0[144:143]!=2'b00));
  assign ensig_cgo_mx0 = nor_cse & (~ (hit_in_crt_sva_171_0[142])) & readHit_sva
      & (or_dcpl_32 | (fsm_output[14]));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_mux_1_cse
      = MUX_s_1_2_2(z_out_21_2, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_acc_1_2_svs_cse,
      z_out_1_33);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_else_if_mux_1_cse
      = MUX_s_1_2_2(z_out_21_2, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_1_2_svs_cse,
      z_out_1_33);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_else_if_mux_1_cse
      & (~ z_out_1_33);
  assign lambertianScatter_run_land_lpi_1_dfm_mx1w0 = (z_out_4[28]) & ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_0;
  assign lambertianScatter_run_if_lambertianScatter_run_if_and_1_nl = (z_out_4[28])
      & lambertianScatter_run_land_1_lpi_1_dfm;
  assign lambertianScatter_run_land_1_lpi_1_dfm_mx2 = MUX_s_1_2_2((lambertianScatter_run_if_lambertianScatter_run_if_and_1_nl),
      lambertianScatter_run_land_1_lpi_1_dfm, or_dcpl_30);
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({(~ reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg)
      , (~ reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg)})
      + 65'b00000000000000000000000000000000000000000000000000000000000000001;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl[64:0];
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_lpi_1_dfm_64_0_mx0
      = MUX_v_65_2_2(({reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg}),
      (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_1_acc_nl),
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1
      = ~(MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), 2'b11, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_else_if_mux_1_cse));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0
      = MUX_v_2_2_2(({{1{z_out_21_2}}, z_out_21_2}), 2'b01, z_out_1_33);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_mux_1_cse
      & (~ z_out_1_33);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1
      = ~(MUX_v_3_2_2(({{2{z_out_1_33}}, z_out_1_33}), 3'b111, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_mux_1_cse));
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva
      + 6'b000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3[5:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva
      + 6'b000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2[5:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1
      = reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg
      + 6'b000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1[5:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2
      = ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva
      + 6'b000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2[5:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl
      = conv_u2s_6_7(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2)
      + 7'b1011011;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl[6:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl
      = conv_u2s_6_7(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_i_5_0_sva_1_mx0w1)
      + 7'b1011011;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl[6:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl
      = conv_u2s_6_7(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2)
      + 7'b1011011;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl[6:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl
      = conv_u2s_6_7(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3)
      + 7'b1011011;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl[6:0];
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_tmp
      = (~((readslicef_7_1_6((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl)))
      | (readslicef_7_1_6((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_acc_nl)))))
      & (~((readslicef_7_1_6((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_acc_nl)))
      | (readslicef_7_1_6((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_acc_nl)))));
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6
      = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0})
      + conv_u2s_42_45(ac_math_atan_pi_2mi_return_69_28_sva);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6[44:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6
      = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0})
      + conv_u2s_42_45(ac_math_atan_pi_2mi_return_1_69_28_sva);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6[44:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6
      = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0})
      + conv_u2s_42_45(ac_math_atan_pi_2mi_return_2_69_28_sva);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6[44:0];
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6
      = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0})
      + conv_u2s_42_45(ac_math_atan_pi_2mi_return_3_69_28_sva);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6[44:0];
  assign and_dcpl_5 = nor_cse & (~ (hit_in_crt_sva_171_0[142]));
  assign and_dcpl_18 = readHit_sva & (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_tmp);
  assign or_dcpl_29 = (hit_in_crt_sva_171_0[144:143]!=2'b00);
  assign or_dcpl_30 = or_dcpl_29 | (hit_in_crt_sva_171_0[142]) | (~ readHit_sva);
  assign or_dcpl_32 = (fsm_output[16:15]!=2'b00);
  assign or_dcpl_35 = or_dcpl_29 | (hit_in_crt_sva_171_0[142]);
  assign or_dcpl_44 = (fsm_output[10]) | (fsm_output[3]);
  assign or_dcpl_45 = or_dcpl_44 | (fsm_output[2]);
  assign and_dcpl_58 = ~((fsm_output[17]) | (fsm_output[15]));
  assign and_dcpl_62 = ~((~ nor_31_cse) | (fsm_output[1]) | (fsm_output[19]) | (fsm_output[18]));
  assign or_dcpl_73 = (fsm_output[16]) | (fsm_output[14]);
  assign or_tmp_44 = (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1)
      & (fsm_output[19]);
  assign or_tmp_54 = (~(readHit_sva & else_unequal_tmp)) & (fsm_output[14]);
  assign or_tmp_78 = readHit_sva & (fsm_output[14]);
  assign or_tmp_111 = readHit_sva & (~ else_unequal_tmp) & (fsm_output[14]);
  assign and_352_cse = ((~ readHit_sva) | else_unequal_tmp) & (fsm_output[14]);
  assign or_tmp_208 = or_dcpl_45 | (fsm_output[4]) | (fsm_output[12]);
  assign or_tmp_400 = (fsm_output[18]) | (fsm_output[17]) | (fsm_output[15]) | or_dcpl_73;
  assign or_tmp_407 = (fsm_output[13:11]!=3'b000);
  assign or_tmp_516 = (fsm_output[10]) | (fsm_output[12]);
  assign or_tmp_659 = ~((fsm_output[13:12]!=2'b00));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs_mx0c2
      = (~ readHit_sva) & (fsm_output[14]);
  assign xor_cse = lambertianScatter_state2_10_sva ^ lambertianScatter_state2_23_sva
      ^ lambertianScatter_state2_6_sva ^ lambertianScatter_state2_11_sva;
  assign rand_unit_random2_run_x3_11_sva_mx0w0 = lambertianScatter_state2_28_sva
      ^ lambertianScatter_state2_15_sva ^ xor_cse;
  assign rand_unit_random2_run_x2_1_sva_mx0w0 = lambertianScatter_state2_1_sva ^
      lambertianScatter_state2_18_sva ^ lambertianScatter_state2_5_sva;
  assign xor_cse_1 = lambertianScatter_state2_9_sva ^ lambertianScatter_state2_22_sva
      ^ lambertianScatter_state2_5_sva ^ lambertianScatter_state2_10_sva;
  assign rand_unit_random2_run_x3_10_sva_mx0w0 = lambertianScatter_state2_27_sva
      ^ lambertianScatter_state2_14_sva ^ xor_cse_1;
  assign rand_unit_random2_run_x2_0_sva_mx0w0 = lambertianScatter_state2_0_sva ^
      lambertianScatter_state2_17_sva ^ lambertianScatter_state2_4_sva;
  assign rand_unit_random2_run_x2_4_sva_mx0w0 = lambertianScatter_state2_4_sva ^
      lambertianScatter_state2_21_sva ^ lambertianScatter_state2_8_sva;
  assign rand_unit_random2_run_x2_3_sva_mx0w0 = lambertianScatter_state2_3_sva ^
      lambertianScatter_state2_20_sva ^ lambertianScatter_state2_7_sva;
  assign rand_unit_random2_run_x2_2_sva_mx0w0 = lambertianScatter_state2_2_sva ^
      lambertianScatter_state2_19_sva ^ lambertianScatter_state2_6_sva;
  assign xor_cse_2 = lambertianScatter_state2_12_sva ^ lambertianScatter_state2_17_sva
      ^ lambertianScatter_state2_4_sva ^ lambertianScatter_state2_29_sva;
  assign rand_unit_random2_run_x3_17_sva_mx0w0 = lambertianScatter_state2_16_sva
      ^ xor_cse_2;
  assign xor_cse_3 = lambertianScatter_state2_15_sva ^ lambertianScatter_state2_28_sva
      ^ lambertianScatter_state2_23_sva;
  assign rand_unit_random2_run_x3_28_sva_mx0w0 = lambertianScatter_state2_10_sva
      ^ xor_cse_3;
  assign xor_cse_4 = lambertianScatter_state2_8_sva ^ lambertianScatter_state2_21_sva
      ^ lambertianScatter_state2_26_sva ^ lambertianScatter_state2_9_sva;
  assign rand_unit_random2_run_x3_9_sva_mx0w0 = lambertianScatter_state2_13_sva ^
      lambertianScatter_state2_4_sva ^ xor_cse_4;
  assign xor_cse_5 = lambertianScatter_state2_4_sva ^ lambertianScatter_state2_9_sva
      ^ lambertianScatter_state2_22_sva ^ lambertianScatter_state2_5_sva;
  assign rand_unit_random2_run_x3_5_sva_mx0w0 = lambertianScatter_state2_0_sva ^
      lambertianScatter_state2_17_sva ^ xor_cse_5;
  assign xor_cse_6 = lambertianScatter_state2_12_sva ^ lambertianScatter_state2_7_sva
      ^ lambertianScatter_state2_25_sva ^ lambertianScatter_state2_8_sva;
  assign rand_unit_random2_run_x3_8_sva_mx0w0 = lambertianScatter_state2_3_sva ^
      lambertianScatter_state2_20_sva ^ xor_cse_6;
  assign xor_cse_7 = lambertianScatter_state2_18_sva ^ lambertianScatter_state2_1_sva
      ^ lambertianScatter_state2_6_sva ^ lambertianScatter_state2_23_sva;
  assign rand_unit_random2_run_x3_6_sva_mx0w0 = lambertianScatter_state2_10_sva ^
      lambertianScatter_state2_5_sva ^ xor_cse_7;
  assign xor_cse_8 = lambertianScatter_state2_11_sva ^ lambertianScatter_state2_24_sva
      ^ lambertianScatter_state2_7_sva ^ lambertianScatter_state2_2_sva;
  assign rand_unit_random2_run_x3_7_sva_mx0w0 = lambertianScatter_state2_19_sva ^
      lambertianScatter_state2_6_sva ^ xor_cse_8;
  assign xor_cse_9 = lambertianScatter_state2_12_sva ^ lambertianScatter_state2_25_sva
      ^ lambertianScatter_state2_30_sva;
  assign rand_unit_random2_run_x3_30_sva_mx0w0 = lambertianScatter_state2_17_sva
      ^ xor_cse_9;
  assign xor_cse_10 = lambertianScatter_state2_14_sva ^ lambertianScatter_state2_27_sva
      ^ lambertianScatter_state2_15_sva ^ lambertianScatter_state2_2_sva;
  assign rand_unit_random2_run_x3_15_sva_mx0w0 = lambertianScatter_state2_10_sva
      ^ xor_cse_10;
  assign xor_cse_11 = lambertianScatter_state2_11_sva ^ lambertianScatter_state2_16_sva
      ^ lambertianScatter_state2_29_sva ^ lambertianScatter_state2_24_sva;
  assign xor_cse_12 = lambertianScatter_state2_13_sva ^ lambertianScatter_state2_26_sva
      ^ lambertianScatter_state2_9_sva ^ lambertianScatter_state2_14_sva;
  assign xor_cse_13 = lambertianScatter_state2_18_sva ^ lambertianScatter_state2_1_sva
      ^ lambertianScatter_state2_31_sva;
  assign rand_unit_random2_run_x3_14_sva_mx0w0 = xor_cse_12 ^ xor_cse_13;
  assign xor_cse_14 = lambertianScatter_state2_22_sva ^ lambertianScatter_state2_9_sva
      ^ lambertianScatter_state2_27_sva;
  assign rand_unit_random2_run_x3_27_sva_mx0w0 = lambertianScatter_state2_14_sva
      ^ xor_cse_14;
  assign xor_cse_15 = lambertianScatter_state2_17_sva ^ lambertianScatter_state2_0_sva
      ^ lambertianScatter_state2_13_sva ^ lambertianScatter_state2_30_sva;
  assign xor_cse_16 = lambertianScatter_state2_8_sva ^ lambertianScatter_state2_25_sva
      ^ lambertianScatter_state2_12_sva;
  assign rand_unit_random2_run_x3_13_sva_mx0w0 = xor_cse_15 ^ xor_cse_16;
  assign rand_unit_random2_run_x3_12_sva_mx0w0 = lambertianScatter_state2_12_sva
      ^ lambertianScatter_state2_7_sva ^ xor_cse_11;
  assign xor_cse_17 = lambertianScatter_state2_8_sva ^ lambertianScatter_state2_21_sva
      ^ lambertianScatter_state2_26_sva;
  assign rand_unit_random2_run_x3_26_sva_mx0w0 = lambertianScatter_state2_13_sva
      ^ xor_cse_17;
  assign xor_cse_18 = lambertianScatter_state2_20_sva ^ lambertianScatter_state2_7_sva
      ^ lambertianScatter_state2_25_sva;
  assign rand_unit_random2_run_x3_25_sva_mx0w0 = lambertianScatter_state2_12_sva
      ^ xor_cse_18;
  assign rand_unit_random2_run_x3_24_sva_mx0w0 = lambertianScatter_state2_24_sva
      ^ lambertianScatter_state2_11_sva ^ lambertianScatter_state2_19_sva ^ lambertianScatter_state2_6_sva;
  assign rand_unit_random2_run_x3_23_sva_mx0w0 = lambertianScatter_state2_23_sva
      ^ lambertianScatter_state2_10_sva ^ lambertianScatter_state2_18_sva ^ lambertianScatter_state2_5_sva;
  assign xor_cse_19 = lambertianScatter_state2_15_sva ^ lambertianScatter_state2_28_sva
      ^ lambertianScatter_state2_16_sva ^ lambertianScatter_state2_3_sva;
  assign rand_unit_random2_run_x3_16_sva_mx0w0 = lambertianScatter_state2_11_sva
      ^ xor_cse_19;
  assign rand_unit_random2_run_x3_22_sva_mx0w0 = lambertianScatter_state2_22_sva
      ^ lambertianScatter_state2_9_sva ^ lambertianScatter_state2_17_sva ^ lambertianScatter_state2_4_sva;
  assign rand_unit_random2_run_x3_18_sva_mx0w0 = lambertianScatter_state2_18_sva
      ^ lambertianScatter_state2_5_sva ^ xor_cse_15;
  assign rand_unit_random2_run_x3_21_sva_mx0w0 = lambertianScatter_state2_21_sva
      ^ lambertianScatter_state2_8_sva ^ lambertianScatter_state2_16_sva ^ lambertianScatter_state2_3_sva;
  assign xor_cse_20 = lambertianScatter_state2_18_sva ^ lambertianScatter_state2_31_sva
      ^ lambertianScatter_state2_1_sva ^ lambertianScatter_state2_19_sva;
  assign rand_unit_random2_run_x3_19_sva_mx0w0 = lambertianScatter_state2_6_sva ^
      lambertianScatter_state2_14_sva ^ xor_cse_20;
  assign rand_unit_random2_run_x3_20_sva_mx0w0 = lambertianScatter_state2_20_sva
      ^ lambertianScatter_state2_7_sva ^ lambertianScatter_state2_15_sva ^ lambertianScatter_state2_2_sva;
  assign rand_unit_random2_run_x3_xor_26_tmp = lambertianScatter_state2_26_sva ^
      lambertianScatter_state2_31_sva ^ lambertianScatter_state2_18_sva ^ lambertianScatter_state2_13_sva;
  assign xor_cse_21 = lambertianScatter_state1_sva_5 ^ lambertianScatter_state1_sva_22
      ^ lambertianScatter_state1_sva_9;
  assign xor_cse_22 = lambertianScatter_state1_sva_12 ^ lambertianScatter_state1_sva_25
      ^ lambertianScatter_state1_sva_20 ^ lambertianScatter_state1_sva_7;
  assign xor_cse_23 = lambertianScatter_state1_sva_10 ^ lambertianScatter_state1_sva_23
      ^ lambertianScatter_state1_sva_6;
  assign xor_cse_24 = lambertianScatter_state1_sva_11 ^ lambertianScatter_state1_sva_24
      ^ lambertianScatter_state1_sva_7;
  assign xor_cse_25 = lambertianScatter_state1_sva_13 ^ lambertianScatter_state1_sva_26
      ^ lambertianScatter_state1_sva_9;
  assign xor_cse_26 = lambertianScatter_state1_sva_14 ^ lambertianScatter_state1_sva_27
      ^ lambertianScatter_state1_sva_10;
  assign xor_cse_27 = lambertianScatter_state1_sva_15 ^ lambertianScatter_state1_sva_28
      ^ lambertianScatter_state1_sva_11;
  assign xor_cse_28 = lambertianScatter_state1_sva_18 ^ lambertianScatter_state1_sva_31
      ^ lambertianScatter_state1_sva_14;
  assign xor_cse_29 = lambertianScatter_state1_sva_16 ^ lambertianScatter_state1_sva_29
      ^ lambertianScatter_state1_sva_12;
  assign xor_cse_30 = lambertianScatter_state1_sva_17 ^ lambertianScatter_state1_sva_0
      ^ lambertianScatter_state1_sva_13 ^ lambertianScatter_state1_sva_30;
  assign lambertianScatter_rand_unit_run_xs_mul_cmp_a = MUX_v_36_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva[42:7]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0,
      fsm_output[15]);
  assign lambertianScatter_rand_unit_run_xs_mul_cmp_b = MUX_v_36_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0,
      fsm_output[15]);
  assign or_tmp_1118 = (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1)
      & (fsm_output[8]);
  assign or_tmp_1119 = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
      & (fsm_output[8]);
  assign and_dcpl_110 = ((fsm_output[7]) | (fsm_output[5]) | (fsm_output[9])) & scatter_wen;
  assign or_1202_ssc = (fsm_output[19:17]!=3'b000);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_cse
      = rand_unit_random1_run_x3_sva_31 | (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_1_cse
      = rand_unit_random1_run_x3_sva_30 | (fsm_output[13]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      ray_out_rsci_idat_41_21 <= 21'b000000000000000000000;
      ray_out_rsci_idat_62_42 <= 21'b000000000000000000000;
      ray_out_rsci_idat_96_63 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_130_97 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_164_131 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_165 <= 1'b0;
    end
    else if ( ray_out_and_cse ) begin
      ray_out_rsci_idat_20_0 <= color_out_r_sva_1_20_0;
      ray_out_rsci_idat_41_21 <= lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0;
      ray_out_rsci_idat_62_42 <= mux_21_itm;
      ray_out_rsci_idat_96_63 <= MUX_v_34_2_2((signext_34_26(lambertianScatter_run_mux_nl)),
          (ray_in_crt_sva[96:63]), or_tmp_44);
      ray_out_rsci_idat_130_97 <= MUX_v_34_2_2((signext_34_26(lambertianScatter_run_mux_1_nl)),
          (ray_in_crt_sva[130:97]), or_tmp_44);
      ray_out_rsci_idat_164_131 <= MUX_v_34_2_2((signext_34_26(lambertianScatter_run_mux_2_nl)),
          (ray_in_crt_sva[164:131]), or_tmp_44);
      ray_out_rsci_idat_165 <= ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_out_rsci_idat_26_0 <= 27'b000000000000000000000000000;
      accumalated_color_out_rsci_idat_53_27 <= 27'b000000000000000000000000000;
      accumalated_color_out_rsci_idat_80_54 <= 27'b000000000000000000000000000;
      attenuation_chan_out_rsci_idat_26_21 <= 6'b000000;
      attenuation_chan_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      attenuation_chan_out_rsci_idat_53_27 <= 27'b000000000000000000000000000;
      attenuation_chan_out_rsci_idat_80 <= 1'b0;
      attenuation_chan_out_rsci_idat_79_54 <= 26'b00000000000000000000000000;
    end
    else if ( accumalated_color_out_and_cse ) begin
      accumalated_color_out_rsci_idat_26_0 <= MUX_v_27_2_2(({color_out_r_sva_1_26_21
          , color_out_r_sva_1_20_0}), (accumalated_color_chan_in_crt_sva[26:0]),
          or_tmp_54);
      accumalated_color_out_rsci_idat_53_27 <= MUX_v_27_2_2(({color_out_g_sva_1_26
          , color_out_g_sva_1_25_0}), (accumalated_color_chan_in_crt_sva[53:27]),
          or_tmp_54);
      accumalated_color_out_rsci_idat_80_54 <= MUX_v_27_2_2(lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0,
          (accumalated_color_chan_in_crt_sva[80:54]), or_tmp_54);
      attenuation_chan_out_rsci_idat_26_21 <= color_out_r_sva_1_26_21 & (signext_6_1(~
          else_unequal_tmp)) & ({{5{readHit_sva}}, readHit_sva});
      attenuation_chan_out_rsci_idat_20_0 <= color_out_r_sva_1_20_0 & (signext_21_1(~
          else_unequal_tmp)) & ({{20{readHit_sva}}, readHit_sva});
      attenuation_chan_out_rsci_idat_53_27 <= lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0
          & (signext_27_1(~ else_unequal_tmp)) & ({{26{readHit_sva}}, readHit_sva});
      attenuation_chan_out_rsci_idat_80 <= color_out_g_sva_1_26 & (~ else_unequal_tmp)
          & readHit_sva;
      attenuation_chan_out_rsci_idat_79_54 <= color_out_g_sva_1_25_0 & (signext_26_1(~
          else_unequal_tmp)) & ({{25{readHit_sva}}, readHit_sva});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ensig_cgo <= 1'b0;
      reg_ray_out_rsci_ivld_scatter_psct_cse <= 1'b0;
      reg_accumalated_color_out_rsci_ivld_scatter_psct_cse <= 1'b0;
      reg_isHit_rsci_irdy_scatter_psct_cse <= 1'b0;
      else_if_mul_cmp_b <= 27'b000000000000000000000000000;
      else_if_mul_cmp_a <= 27'b000000000000000000000000000;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16
          <= 1'b0;
      hit_in_crt_sva_198_172 <= 27'b000000000000000000000000000;
      attenuation_chan_in_crt_sva_53_27 <= 27'b000000000000000000000000000;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva <= 69'b000000000000000000000000000000000000000000000000000000000000000000000;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_7_4
          <= 4'b0000;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_sva
          <= 69'b000000000000000000000000000000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0
          <= 36'b000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0
          <= 36'b000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs
          <= 1'b0;
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd
          <= 2'b00;
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1
          <= 26'b00000000000000000000000000;
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_3
          <= 7'b0000000;
    end
    else if ( scatter_wen ) begin
      ensig_cgo <= ensig_cgo_mx0;
      reg_ray_out_rsci_ivld_scatter_psct_cse <= fsm_output[19];
      reg_accumalated_color_out_rsci_ivld_scatter_psct_cse <= fsm_output[14];
      reg_isHit_rsci_irdy_scatter_psct_cse <= ~ nor_31_cse;
      else_if_mul_cmp_b <= MUX1HOT_v_27_3_2((hit_in_rsci_idat_mxwt[225:199]), hit_in_crt_sva_198_172,
          (hit_in_crt_sva_171_0[171:145]), {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[3])});
      else_if_mul_cmp_a <= MUX1HOT_v_27_3_2((attenuation_chan_in_rsci_idat_mxwt[80:54]),
          attenuation_chan_in_crt_sva_53_27, attenuation_chan_in_crt_sva_26_0, {(fsm_output[1])
          , (fsm_output[2]) , (fsm_output[3])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_4_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_8_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_17_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_41_nl)
          & (~ (fsm_output[11]));
      hit_in_crt_sva_198_172 <= hit_in_rsci_idat_mxwt[198:172];
      attenuation_chan_in_crt_sva_53_27 <= attenuation_chan_in_rsci_idat_mxwt[53:27];
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva <= nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva[68:0];
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_7_4
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_rgt[7:4];
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_sva
          <= z_out_19;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux1h_89_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_33_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_32_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_7_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_2_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0
          <= MUX_v_36_2_2(36'b000000000000000000000000000000000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_16_nl),
          (not_319_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_6_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_5_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_4_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_3_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_2_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_1_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11
          <= (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0
          <= MUX_v_36_2_2(36'b000000000000000000000000000000000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_15_nl),
          (not_306_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_10_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_6_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11
          <= (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl)
          & (~ (fsm_output[11]));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva
          <= MUX_v_43_2_2((z_out_19[42:0]), ({(z_out_12[42:7]) , 7'b0000000}), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm
          <= ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_tmp;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs
          <= MUX_s_1_2_2((z_out_8[45]), lambertianScatter_run_land_lpi_1_dfm_mx1w0,
          fsm_output[18]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs
          <= z_out_9[45];
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd
          <= operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm[42:41];
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1
          <= MUX_v_26_2_2((operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm[40:15]),
          (z_out_10[40:15]), fsm_output[13]);
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_3
          <= operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm[6:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_acc_1_2_svs_cse
          <= 1'b0;
    end
    else if ( scatter_wen & (~((~ (fsm_output[11])) | or_dcpl_35 | (~ readHit_sva)
        | z_out_1_33)) ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_else_if_acc_1_2_svs_cse
          <= z_out_21_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_state2_0_sva <= 1'b0;
      lambertianScatter_state2_1_sva <= 1'b0;
      lambertianScatter_state2_2_sva <= 1'b0;
      lambertianScatter_state2_3_sva <= 1'b0;
      lambertianScatter_state2_4_sva <= 1'b1;
      lambertianScatter_state2_5_sva <= 1'b0;
      lambertianScatter_state2_6_sva <= 1'b0;
      lambertianScatter_state2_7_sva <= 1'b1;
      lambertianScatter_state2_8_sva <= 1'b0;
      lambertianScatter_state2_9_sva <= 1'b0;
      lambertianScatter_state2_10_sva <= 1'b1;
      lambertianScatter_state2_11_sva <= 1'b1;
      lambertianScatter_state2_12_sva <= 1'b0;
      lambertianScatter_state2_13_sva <= 1'b1;
      lambertianScatter_state2_14_sva <= 1'b1;
      lambertianScatter_state2_16_sva <= 1'b0;
      lambertianScatter_state2_15_sva <= 1'b1;
      lambertianScatter_state2_31_sva <= 1'b0;
      lambertianScatter_state2_18_sva <= 1'b1;
      lambertianScatter_state2_30_sva <= 1'b0;
      lambertianScatter_state2_17_sva <= 1'b1;
      lambertianScatter_state2_29_sva <= 1'b0;
      lambertianScatter_state2_28_sva <= 1'b0;
      lambertianScatter_state2_27_sva <= 1'b0;
      lambertianScatter_state2_26_sva <= 1'b0;
      lambertianScatter_state2_25_sva <= 1'b1;
      lambertianScatter_state2_24_sva <= 1'b0;
      lambertianScatter_state2_23_sva <= 1'b0;
      lambertianScatter_state2_22_sva <= 1'b1;
      lambertianScatter_state2_21_sva <= 1'b0;
      lambertianScatter_state2_20_sva <= 1'b1;
      lambertianScatter_state2_19_sva <= 1'b0;
    end
    else if ( lambertianScatter_state2_and_32_cse ) begin
      lambertianScatter_state2_0_sva <= lambertianScatter_state1_sva_0;
      lambertianScatter_state2_1_sva <= lambertianScatter_state1_sva_1;
      lambertianScatter_state2_2_sva <= lambertianScatter_state1_sva_10;
      lambertianScatter_state2_3_sva <= lambertianScatter_state1_sva_11;
      lambertianScatter_state2_4_sva <= lambertianScatter_state1_sva_12;
      lambertianScatter_state2_5_sva <= lambertianScatter_state1_sva_4;
      lambertianScatter_state2_6_sva <= lambertianScatter_state1_sva_5;
      lambertianScatter_state2_7_sva <= lambertianScatter_state1_sva_6;
      lambertianScatter_state2_8_sva <= lambertianScatter_state1_sva_7;
      lambertianScatter_state2_9_sva <= lambertianScatter_state1_sva_8;
      lambertianScatter_state2_10_sva <= lambertianScatter_state1_sva_13;
      lambertianScatter_state2_11_sva <= lambertianScatter_state1_sva_14;
      lambertianScatter_state2_12_sva <= lambertianScatter_state1_sva_15;
      lambertianScatter_state2_13_sva <= lambertianScatter_state1_sva_16;
      lambertianScatter_state2_14_sva <= lambertianScatter_state1_sva_17;
      lambertianScatter_state2_16_sva <= lambertianScatter_state1_sva_19;
      lambertianScatter_state2_15_sva <= lambertianScatter_state1_sva_18;
      lambertianScatter_state2_31_sva <= rand_unit_random2_run_x3_31_sva;
      lambertianScatter_state2_18_sva <= lambertianScatter_state1_sva_20;
      lambertianScatter_state2_30_sva <= lambertianScatter_state1_sva_31;
      lambertianScatter_state2_17_sva <= lambertianScatter_state1_sva_2;
      lambertianScatter_state2_29_sva <= lambertianScatter_state1_sva_30;
      lambertianScatter_state2_28_sva <= lambertianScatter_state1_sva_3;
      lambertianScatter_state2_27_sva <= lambertianScatter_state1_sva_29;
      lambertianScatter_state2_26_sva <= lambertianScatter_state1_sva_28;
      lambertianScatter_state2_25_sva <= lambertianScatter_state1_sva_27;
      lambertianScatter_state2_24_sva <= lambertianScatter_state1_sva_26;
      lambertianScatter_state2_23_sva <= lambertianScatter_state1_sva_25;
      lambertianScatter_state2_22_sva <= lambertianScatter_state1_sva_24;
      lambertianScatter_state2_21_sva <= lambertianScatter_state1_sva_23;
      lambertianScatter_state2_20_sva <= lambertianScatter_state1_sva_22;
      lambertianScatter_state2_19_sva <= lambertianScatter_state1_sva_21;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_state1_sva_14 <= 1'b0;
      lambertianScatter_state1_sva_1 <= 1'b0;
      lambertianScatter_state1_sva_13 <= 1'b1;
      lambertianScatter_state1_sva_0 <= 1'b1;
      lambertianScatter_state1_sva_12 <= 1'b1;
      lambertianScatter_state1_sva_11 <= 1'b1;
      lambertianScatter_state1_sva_10 <= 1'b1;
      lambertianScatter_state1_sva_2 <= 1'b1;
      lambertianScatter_state1_sva_3 <= 1'b1;
      lambertianScatter_state1_sva_8 <= 1'b0;
      lambertianScatter_state1_sva_4 <= 1'b0;
      lambertianScatter_state1_sva_7 <= 1'b0;
      lambertianScatter_state1_sva_5 <= 1'b0;
      lambertianScatter_state1_sva_6 <= 1'b0;
      lambertianScatter_state1_sva_31 <= 1'b0;
      lambertianScatter_state1_sva_18 <= 1'b1;
      lambertianScatter_state1_sva_30 <= 1'b0;
      lambertianScatter_state1_sva_17 <= 1'b0;
      lambertianScatter_state1_sva_29 <= 1'b0;
      lambertianScatter_state1_sva_16 <= 1'b1;
      lambertianScatter_state1_sva_15 <= 1'b1;
      lambertianScatter_state1_sva_28 <= 1'b0;
      lambertianScatter_state1_sva_27 <= 1'b0;
      lambertianScatter_state1_sva_26 <= 1'b0;
      lambertianScatter_state1_sva_25 <= 1'b0;
      lambertianScatter_state1_sva_19 <= 1'b0;
      lambertianScatter_state1_sva_24 <= 1'b0;
      lambertianScatter_state1_sva_20 <= 1'b0;
      lambertianScatter_state1_sva_23 <= 1'b0;
      lambertianScatter_state1_sva_21 <= 1'b0;
      lambertianScatter_state1_sva_22 <= 1'b0;
    end
    else if ( lambertianScatter_state1_and_cse ) begin
      lambertianScatter_state1_sva_14 <= MUX_s_1_2_2(rand_unit_random2_run_x3_11_sva_mx0w0,
          rand_unit_random1_run_x3_sva_14, or_tmp_111);
      lambertianScatter_state1_sva_1 <= MUX_s_1_2_2(rand_unit_random2_run_x2_1_sva_mx0w0,
          rand_unit_random1_run_x2_12_0_sva_1, or_tmp_111);
      lambertianScatter_state1_sva_13 <= MUX_s_1_2_2(rand_unit_random2_run_x3_10_sva_mx0w0,
          rand_unit_random1_run_x3_sva_13, or_tmp_111);
      lambertianScatter_state1_sva_0 <= MUX_s_1_2_2(rand_unit_random2_run_x2_0_sva_mx0w0,
          rand_unit_random1_run_x2_12_0_sva_0, or_tmp_111);
      lambertianScatter_state1_sva_12 <= MUX_s_1_2_2(rand_unit_random2_run_x2_4_sva_mx0w0,
          rand_unit_random1_run_x3_sva_12, or_tmp_111);
      lambertianScatter_state1_sva_11 <= MUX_s_1_2_2(rand_unit_random2_run_x2_3_sva_mx0w0,
          rand_unit_random1_run_x3_sva_11, or_tmp_111);
      lambertianScatter_state1_sva_10 <= MUX_s_1_2_2(rand_unit_random2_run_x2_2_sva_mx0w0,
          rand_unit_random1_run_x3_sva_10, or_tmp_111);
      lambertianScatter_state1_sva_2 <= MUX_s_1_2_2(rand_unit_random2_run_x3_17_sva_mx0w0,
          rand_unit_random1_run_x2_12_0_sva_2, or_tmp_111);
      lambertianScatter_state1_sva_3 <= MUX_s_1_2_2(rand_unit_random2_run_x3_28_sva_mx0w0,
          rand_unit_random1_run_x2_12_0_sva_3, or_tmp_111);
      lambertianScatter_state1_sva_8 <= MUX_s_1_2_2(rand_unit_random2_run_x3_9_sva_mx0w0,
          rand_unit_random1_run_x3_sva_8, or_tmp_111);
      lambertianScatter_state1_sva_4 <= MUX_s_1_2_2(rand_unit_random2_run_x3_5_sva_mx0w0,
          rand_unit_random1_run_x2_12_0_sva_4, or_tmp_111);
      lambertianScatter_state1_sva_7 <= MUX_s_1_2_2(rand_unit_random2_run_x3_8_sva_mx0w0,
          rand_unit_random1_run_x3_sva_7, or_tmp_111);
      lambertianScatter_state1_sva_5 <= MUX_s_1_2_2(rand_unit_random2_run_x3_6_sva_mx0w0,
          rand_unit_random1_run_x3_sva_5, or_tmp_111);
      lambertianScatter_state1_sva_6 <= MUX_s_1_2_2(rand_unit_random2_run_x3_7_sva_mx0w0,
          rand_unit_random1_run_x3_sva_6, or_tmp_111);
      lambertianScatter_state1_sva_31 <= MUX_s_1_2_2(rand_unit_random2_run_x3_30_sva_mx0w0,
          rand_unit_random1_run_x3_sva_31, or_tmp_111);
      lambertianScatter_state1_sva_18 <= MUX_s_1_2_2(rand_unit_random2_run_x3_15_sva_mx0w0,
          rand_unit_random1_run_x3_sva_18, or_tmp_111);
      lambertianScatter_state1_sva_30 <= MUX_s_1_2_2(xor_cse_11, rand_unit_random1_run_x3_sva_30,
          or_tmp_111);
      lambertianScatter_state1_sva_17 <= MUX_s_1_2_2(rand_unit_random2_run_x3_14_sva_mx0w0,
          rand_unit_random1_run_x3_sva_17, or_tmp_111);
      lambertianScatter_state1_sva_29 <= MUX_s_1_2_2(rand_unit_random2_run_x3_27_sva_mx0w0,
          rand_unit_random1_run_x3_sva_29, or_tmp_111);
      lambertianScatter_state1_sva_16 <= MUX_s_1_2_2(rand_unit_random2_run_x3_13_sva_mx0w0,
          rand_unit_random1_run_x3_sva_16, or_tmp_111);
      lambertianScatter_state1_sva_15 <= MUX_s_1_2_2(rand_unit_random2_run_x3_12_sva_mx0w0,
          rand_unit_random1_run_x3_sva_15, or_tmp_111);
      lambertianScatter_state1_sva_28 <= MUX_s_1_2_2(rand_unit_random2_run_x3_26_sva_mx0w0,
          rand_unit_random1_run_x3_sva_28, or_tmp_111);
      lambertianScatter_state1_sva_27 <= MUX_s_1_2_2(rand_unit_random2_run_x3_25_sva_mx0w0,
          rand_unit_random1_run_x3_sva_27, or_tmp_111);
      lambertianScatter_state1_sva_26 <= MUX_s_1_2_2(rand_unit_random2_run_x3_24_sva_mx0w0,
          rand_unit_random1_run_x3_sva_26, or_tmp_111);
      lambertianScatter_state1_sva_25 <= MUX_s_1_2_2(rand_unit_random2_run_x3_23_sva_mx0w0,
          rand_unit_random1_run_x3_sva_25, or_tmp_111);
      lambertianScatter_state1_sva_19 <= MUX_s_1_2_2(rand_unit_random2_run_x3_16_sva_mx0w0,
          rand_unit_random1_run_x3_sva_19, or_tmp_111);
      lambertianScatter_state1_sva_24 <= MUX_s_1_2_2(rand_unit_random2_run_x3_22_sva_mx0w0,
          rand_unit_random1_run_x3_sva_24, or_tmp_111);
      lambertianScatter_state1_sva_20 <= MUX_s_1_2_2(rand_unit_random2_run_x3_18_sva_mx0w0,
          rand_unit_random1_run_x3_sva_20, or_tmp_111);
      lambertianScatter_state1_sva_23 <= MUX_s_1_2_2(rand_unit_random2_run_x3_21_sva_mx0w0,
          rand_unit_random1_run_x3_sva_23, or_tmp_111);
      lambertianScatter_state1_sva_21 <= MUX_s_1_2_2(rand_unit_random2_run_x3_19_sva_mx0w0,
          rand_unit_random1_run_x3_sva_21, or_tmp_111);
      lambertianScatter_state1_sva_22 <= MUX_s_1_2_2(rand_unit_random2_run_x3_20_sva_mx0w0,
          rand_unit_random1_run_x3_sva_22, or_tmp_111);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_state1_sva_9 <= 1'b0;
    end
    else if ( scatter_wen & or_tmp_111 ) begin
      lambertianScatter_state1_sva_9 <= rand_unit_random1_run_x3_sva_9;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_1_2_svs_cse
          <= 1'b0;
    end
    else if ( scatter_wen & (~((~ (fsm_output[9])) | or_dcpl_35 | (~ readHit_sva)
        | z_out_1_33)) ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_slc_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_1_2_svs_cse
          <= z_out_21_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12
          <= 1'b0;
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14
          <= 1'b0;
    end
    else if ( ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_45_cse
        ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7
          <= MUX1HOT_s_1_5_2((z_out_3[7]), rand_unit_random2_run_x3_7_sva_mx0w0,
          z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[20]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8
          <= MUX1HOT_s_1_5_2((z_out_3[8]), rand_unit_random2_run_x3_8_sva_mx0w0,
          z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[21]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9
          <= MUX1HOT_s_1_5_2((z_out_3[9]), rand_unit_random2_run_x3_9_sva_mx0w0,
          z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[22]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20
          <= MUX1HOT_s_1_5_2((z_out_3[20]), rand_unit_random2_run_x3_20_sva_mx0w0,
          z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[12]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12
          <= MUX1HOT_s_1_5_2((z_out_3[12]), rand_unit_random2_run_x3_12_sva_mx0w0,
          z_out_1_33, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_0,
          (z_out_14[0]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14
          <= MUX1HOT_s_1_5_2((z_out_3[14]), rand_unit_random2_run_x3_14_sva_mx0w0,
          z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[10]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rand_unit_random2_run_x3_31_sva <= 1'b0;
      rand_unit_random1_run_x3_sva_31 <= 1'b0;
      rand_unit_random1_run_x3_sva_30 <= 1'b0;
      rand_unit_random1_run_x3_sva_29 <= 1'b0;
      rand_unit_random1_run_x3_sva_28 <= 1'b0;
      rand_unit_random1_run_x3_sva_27 <= 1'b0;
      rand_unit_random1_run_x3_sva_26 <= 1'b0;
      rand_unit_random1_run_x3_sva_5 <= 1'b0;
      rand_unit_random1_run_x2_12_0_sva_0 <= 1'b0;
      rand_unit_random1_run_x3_sva_25 <= 1'b0;
      rand_unit_random1_run_x3_sva_6 <= 1'b0;
      rand_unit_random1_run_x2_12_0_sva_1 <= 1'b0;
      rand_unit_random1_run_x3_sva_24 <= 1'b0;
      rand_unit_random1_run_x3_sva_7 <= 1'b0;
      rand_unit_random1_run_x2_12_0_sva_2 <= 1'b0;
      rand_unit_random1_run_x3_sva_23 <= 1'b0;
      rand_unit_random1_run_x3_sva_8 <= 1'b0;
      rand_unit_random1_run_x2_12_0_sva_3 <= 1'b0;
      rand_unit_random1_run_x3_sva_22 <= 1'b0;
      rand_unit_random1_run_x3_sva_9 <= 1'b0;
      rand_unit_random1_run_x2_12_0_sva_4 <= 1'b0;
      rand_unit_random1_run_x3_sva_21 <= 1'b0;
      rand_unit_random1_run_x3_sva_10 <= 1'b0;
      rand_unit_random1_run_x3_sva_20 <= 1'b0;
      rand_unit_random1_run_x3_sva_11 <= 1'b0;
      rand_unit_random1_run_x3_sva_19 <= 1'b0;
      rand_unit_random1_run_x3_sva_12 <= 1'b0;
      rand_unit_random1_run_x3_sva_18 <= 1'b0;
      rand_unit_random1_run_x3_sva_13 <= 1'b0;
      rand_unit_random1_run_x3_sva_17 <= 1'b0;
      rand_unit_random1_run_x3_sva_14 <= 1'b0;
      rand_unit_random1_run_x3_sva_16 <= 1'b0;
      rand_unit_random1_run_x3_sva_15 <= 1'b0;
      accumalated_color_chan_in_crt_sva <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rand_unit_random2_run_x3_and_cse ) begin
      rand_unit_random2_run_x3_31_sva <= rand_unit_random2_run_x3_xor_26_tmp;
      rand_unit_random1_run_x3_sva_31 <= lambertianScatter_state1_sva_31 ^ lambertianScatter_state1_sva_18
          ^ lambertianScatter_state1_sva_26 ^ lambertianScatter_state1_sva_13;
      rand_unit_random1_run_x3_sva_30 <= lambertianScatter_state1_sva_30 ^ lambertianScatter_state1_sva_17
          ^ lambertianScatter_state1_sva_25 ^ lambertianScatter_state1_sva_12;
      rand_unit_random1_run_x3_sva_29 <= lambertianScatter_state1_sva_29 ^ lambertianScatter_state1_sva_16
          ^ lambertianScatter_state1_sva_24 ^ lambertianScatter_state1_sva_11;
      rand_unit_random1_run_x3_sva_28 <= lambertianScatter_state1_sva_28 ^ lambertianScatter_state1_sva_15
          ^ lambertianScatter_state1_sva_23 ^ lambertianScatter_state1_sva_10;
      rand_unit_random1_run_x3_sva_27 <= lambertianScatter_state1_sva_27 ^ lambertianScatter_state1_sva_14
          ^ lambertianScatter_state1_sva_22 ^ lambertianScatter_state1_sva_9;
      rand_unit_random1_run_x3_sva_26 <= lambertianScatter_state1_sva_26 ^ lambertianScatter_state1_sva_13
          ^ lambertianScatter_state1_sva_21 ^ lambertianScatter_state1_sva_8;
      rand_unit_random1_run_x3_sva_5 <= lambertianScatter_state1_sva_0 ^ lambertianScatter_state1_sva_17
          ^ lambertianScatter_state1_sva_4 ^ xor_cse_21;
      rand_unit_random1_run_x2_12_0_sva_0 <= lambertianScatter_state1_sva_0 ^ lambertianScatter_state1_sva_17
          ^ lambertianScatter_state1_sva_4;
      rand_unit_random1_run_x3_sva_25 <= xor_cse_22;
      rand_unit_random1_run_x3_sva_6 <= lambertianScatter_state1_sva_1 ^ lambertianScatter_state1_sva_18
          ^ lambertianScatter_state1_sva_5 ^ xor_cse_23;
      rand_unit_random1_run_x2_12_0_sva_1 <= lambertianScatter_state1_sva_1 ^ lambertianScatter_state1_sva_18
          ^ lambertianScatter_state1_sva_5;
      rand_unit_random1_run_x3_sva_24 <= lambertianScatter_state1_sva_24 ^ lambertianScatter_state1_sva_11
          ^ lambertianScatter_state1_sva_19 ^ lambertianScatter_state1_sva_6;
      rand_unit_random1_run_x3_sva_7 <= lambertianScatter_state1_sva_2 ^ lambertianScatter_state1_sva_19
          ^ lambertianScatter_state1_sva_6 ^ xor_cse_24;
      rand_unit_random1_run_x2_12_0_sva_2 <= lambertianScatter_state1_sva_2 ^ lambertianScatter_state1_sva_19
          ^ lambertianScatter_state1_sva_6;
      rand_unit_random1_run_x3_sva_23 <= lambertianScatter_state1_sva_23 ^ lambertianScatter_state1_sva_10
          ^ lambertianScatter_state1_sva_18 ^ lambertianScatter_state1_sva_5;
      rand_unit_random1_run_x3_sva_8 <= lambertianScatter_state1_sva_8 ^ lambertianScatter_state1_sva_3
          ^ xor_cse_22;
      rand_unit_random1_run_x2_12_0_sva_3 <= lambertianScatter_state1_sva_3 ^ lambertianScatter_state1_sva_20
          ^ lambertianScatter_state1_sva_7;
      rand_unit_random1_run_x3_sva_22 <= lambertianScatter_state1_sva_22 ^ lambertianScatter_state1_sva_9
          ^ lambertianScatter_state1_sva_17 ^ lambertianScatter_state1_sva_4;
      rand_unit_random1_run_x3_sva_9 <= lambertianScatter_state1_sva_4 ^ lambertianScatter_state1_sva_21
          ^ lambertianScatter_state1_sva_8 ^ xor_cse_25;
      rand_unit_random1_run_x2_12_0_sva_4 <= lambertianScatter_state1_sva_4 ^ lambertianScatter_state1_sva_21
          ^ lambertianScatter_state1_sva_8;
      rand_unit_random1_run_x3_sva_21 <= lambertianScatter_state1_sva_21 ^ lambertianScatter_state1_sva_8
          ^ lambertianScatter_state1_sva_16 ^ lambertianScatter_state1_sva_3;
      rand_unit_random1_run_x3_sva_10 <= xor_cse_26 ^ xor_cse_21;
      rand_unit_random1_run_x3_sva_20 <= lambertianScatter_state1_sva_20 ^ lambertianScatter_state1_sva_7
          ^ lambertianScatter_state1_sva_15 ^ lambertianScatter_state1_sva_2;
      rand_unit_random1_run_x3_sva_11 <= xor_cse_23 ^ xor_cse_27;
      rand_unit_random1_run_x3_sva_19 <= lambertianScatter_state1_sva_19 ^ lambertianScatter_state1_sva_6
          ^ lambertianScatter_state1_sva_1 ^ xor_cse_28;
      rand_unit_random1_run_x3_sva_12 <= xor_cse_24 ^ xor_cse_29;
      rand_unit_random1_run_x3_sva_18 <= lambertianScatter_state1_sva_18 ^ lambertianScatter_state1_sva_5
          ^ xor_cse_30;
      rand_unit_random1_run_x3_sva_13 <= lambertianScatter_state1_sva_8 ^ lambertianScatter_state1_sva_25
          ^ lambertianScatter_state1_sva_12 ^ xor_cse_30;
      rand_unit_random1_run_x3_sva_17 <= lambertianScatter_state1_sva_17 ^ lambertianScatter_state1_sva_4
          ^ xor_cse_29;
      rand_unit_random1_run_x3_sva_14 <= lambertianScatter_state1_sva_1 ^ xor_cse_25
          ^ xor_cse_28;
      rand_unit_random1_run_x3_sva_16 <= lambertianScatter_state1_sva_16 ^ lambertianScatter_state1_sva_3
          ^ xor_cse_27;
      rand_unit_random1_run_x3_sva_15 <= lambertianScatter_state1_sva_15 ^ lambertianScatter_state1_sva_2
          ^ xor_cse_26;
      accumalated_color_chan_in_crt_sva <= accumalated_color_chan_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_add_run_acc_4_psp_sva <= 27'b000000000000000000000000000;
    end
    else if ( scatter_wen & (~ or_dcpl_35) & (fsm_output[14]) ) begin
      lambertianScatter_add_run_acc_4_psp_sva <= z_out_15[26:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_run_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( scatter_wen & (~ or_dcpl_30) & (fsm_output[18]) ) begin
      lambertianScatter_run_land_1_lpi_1_dfm <= lambertianScatter_run_land_lpi_1_dfm_mx1w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      else_unequal_tmp <= 1'b0;
      readHit_sva <= 1'b0;
    end
    else if ( else_and_cse ) begin
      else_unequal_tmp <= (hit_in_rsci_idat_mxwt[144:142]!=3'b000);
      readHit_sva <= isHit_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      hit_in_crt_sva_171_0 <= 172'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ((fsm_output[20]) | (fsm_output[0]) | (fsm_output[19]) | (fsm_output[1]))
        & scatter_wen ) begin
      hit_in_crt_sva_171_0 <= hit_in_rsci_idat_mxwt[171:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan_in_crt_sva_26_0 <= 27'b000000000000000000000000000;
    end
    else if ( (~ (fsm_output[2])) & scatter_wen ) begin
      attenuation_chan_in_crt_sva_26_0 <= attenuation_chan_in_rsci_idat_mxwt[26:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_in_crt_sva <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( scatter_wen & (~(nor_31_cse & (~ (fsm_output[1])) & (~ (fsm_output[19]))))
        ) begin
      ray_in_crt_sva <= ray_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14
          <= 2'b00;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_84_cse
        ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11
          <= MUX1HOT_s_1_4_2((z_out_3[1]), rand_unit_random2_run_x2_1_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[11]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12
          <= MUX1HOT_s_1_4_2((z_out_3[10]), rand_unit_random2_run_x3_10_sva_mx0w0,
          z_out_1_33, (z_out_15[12]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13
          <= MUX1HOT_s_1_4_2((z_out_3[11]), rand_unit_random2_run_x3_11_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[13]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16
          <= MUX1HOT_s_1_4_2((z_out_3[13]), rand_unit_random2_run_x3_13_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[16]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19
          <= MUX1HOT_s_1_4_2((z_out_3[15]), rand_unit_random2_run_x3_15_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[19]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23
          <= MUX1HOT_s_1_4_2((z_out_3[17]), rand_unit_random2_run_x3_17_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[23]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24
          <= MUX1HOT_s_1_4_2((z_out_3[18]), rand_unit_random2_run_x3_18_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[24]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25
          <= MUX1HOT_s_1_4_2((z_out_3[19]), rand_unit_random2_run_x3_19_sva_mx0w0,
          z_out_1_33, (z_out_15[25]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26
          <= MUX1HOT_s_1_4_2((z_out_3[2]), rand_unit_random2_run_x2_2_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[26]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30
          <= MUX1HOT_s_1_4_2((z_out_3[21]), rand_unit_random2_run_x3_21_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[30]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33
          <= MUX1HOT_s_1_4_2((z_out_3[23]), rand_unit_random2_run_x3_23_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[33]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36
          <= MUX1HOT_s_1_4_2((z_out_3[25]), rand_unit_random2_run_x3_25_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[36]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37
          <= MUX1HOT_s_1_4_2((z_out_3[26]), rand_unit_random2_run_x3_26_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[37]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38
          <= MUX1HOT_s_1_4_2((z_out_3[27]), rand_unit_random2_run_x3_27_sva_mx0w0,
          z_out_1_33, (z_out_15[38]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5
          <= MUX1HOT_s_1_4_2((z_out_3[29]), xor_cse_11, z_out_1_33, (z_out_15[5]),
          {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6
          <= MUX1HOT_s_1_4_2((z_out_3[3]), rand_unit_random2_run_x2_3_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[6]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7
          <= MUX1HOT_s_1_4_2((z_out_3[4]), rand_unit_random2_run_x2_4_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[7]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8
          <= MUX1HOT_s_1_4_2((z_out_3[5]), rand_unit_random2_run_x3_5_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[8]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9
          <= MUX1HOT_s_1_4_2((z_out_3[6]), rand_unit_random2_run_x3_6_sva_mx0w0,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_15[9]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14
          <= MUX1HOT_v_2_4_2((z_out_3[31:30]), ({1'b0 , rand_unit_random2_run_x3_30_sva_mx0w0}),
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_14[15:14]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[9]) , (fsm_output[13])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm
          <= 1'b0;
    end
    else if ( scatter_wen & (~(or_dcpl_44 | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[7])
        | (fsm_output[11]) | (fsm_output[12]))) ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm
          <= MUX1HOT_s_1_5_2((z_out_3[0]), rand_unit_random2_run_x2_0_sva_mx0w0,
          (readslicef_7_1_6((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl))),
          z_out_1_33, (z_out_15[10]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
          , (fsm_output[6]) , (fsm_output[9]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_out_g_sva_1_26 <= 1'b0;
    end
    else if ( ((fsm_output[15]) | (fsm_output[3]) | (fsm_output[16]) | color_out_g_and_1_cse)
        & scatter_wen ) begin
      color_out_g_sva_1_26 <= color_out_g_mux1h_5_rgt[26];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_out_g_sva_1_25_0 <= 26'b00000000000000000000000000;
    end
    else if ( ((fsm_output[15]) | (fsm_output[3]) | color_out_g_and_1_cse) & scatter_wen
        ) begin
      color_out_g_sva_1_25_0 <= color_out_g_mux1h_5_rgt[25:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_27 <= 1'b0;
    end
    else if ( (~((fsm_output[20]) | (fsm_output[0]) | (fsm_output[19]))) & (~((fsm_output[1])
        | (fsm_output[14]) | (fsm_output[2]))) & scatter_wen ) begin
      lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_27 <= lambertianScatter_run_aelse_1_mux1h_7_rgt[27];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0 <=
          27'b000000000000000000000000000;
    end
    else if ( (color_out_g_and_cse | (fsm_output[3]) | (fsm_output[18]) | (fsm_output[16])
        | (fsm_output[15]) | (fsm_output[17])) & scatter_wen ) begin
      lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0 <=
          lambertianScatter_run_aelse_1_mux1h_7_rgt[26:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_out_r_sva_1_26_21 <= 6'b000000;
    end
    else if ( ((fsm_output[15]) | (fsm_output[16]) | (fsm_output[18]) | (fsm_output[17])
        | (fsm_output[14]) | (fsm_output[5])) & scatter_wen ) begin
      color_out_r_sva_1_26_21 <= color_out_r_mux1h_3_rgt[26:21];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      color_out_r_sva_1_20_0 <= 21'b000000000000000000000;
    end
    else if ( ((fsm_output[14]) | (fsm_output[5])) & scatter_wen ) begin
      color_out_r_sva_1_20_0 <= color_out_r_mux1h_3_rgt[20:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65
          <= 1'b0;
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg
          <= 32'b00000000000000000000000000000000;
    end
    else if ( and_dcpl_110 ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_rgt[65];
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_2_reg
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_rgt[31:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg
          <= 33'b000000000000000000000000000000000;
    end
    else if ( ((fsm_output[7]) | (fsm_output[5]) | ((fsm_output[9]) & ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65))
        & scatter_wen ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_1_reg
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_rgt[64:32];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg
          <= 1'b0;
    end
    else if ( ((fsm_output[11]) | (fsm_output[12]) | (fsm_output[8]) | (fsm_output[5])
        | (fsm_output[13])) & scatter_wen ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_rgt[6];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg
          <= 6'b000000;
    end
    else if ( ((fsm_output[11]) | (fsm_output[12]) | (fsm_output[8]) | (fsm_output[5]))
        & scatter_wen ) begin
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_and_rgt[5:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva <=
          69'b000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( scatter_wen & ((fsm_output[7]) | (fsm_output[8]) | (fsm_output[5]))
        ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva <=
          MUX1HOT_v_69_3_2(69'b001000000000000000000000000000000000000000000000000000000000000000000,
          (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl),
          (z_out_5[68:0]), {(fsm_output[5]) , (fsm_output[7]) , (fsm_output[8])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva <=
          69'b000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( scatter_wen & ((fsm_output[8]) | (fsm_output[5])) ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva <=
          MUX_v_69_2_2(({2'b00 , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11
          , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm
          , 35'b00000000000000000000000000000000000}), (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl),
          fsm_output[8]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm
          <= 69'b000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( (~((fsm_output[6]) | (fsm_output[8]))) & scatter_wen ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm
          <= MUX_v_69_2_2(69'b000000000000000000000000000000000000000000000000000000000000000000000,
          (z_out_5[68:0]), (not_341_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
          <= 1'b0;
    end
    else if ( scatter_wen & ((fsm_output[9]) | (fsm_output[6]) | (fsm_output[8])
        | (fsm_output[12]) | (fsm_output[14])) ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
          <= MUX1HOT_s_1_5_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_or_nl),
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_sva_65,
          (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_nor_nl),
          (z_out_6[45]), and_8_cse, {(fsm_output[6]) , (fsm_output[8]) , (fsm_output[9])
          , (fsm_output[12]) , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_x2_acos_pi_2mi_64_return_sva <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_x_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_theta_d_and_cse
        ) begin
      ac_math_x2_acos_pi_2mi_64_return_sva <= MUX_v_64_66_2(64'b1000000000000000000000000000000000000000000000000000000000000000,
          64'b0100101110010000000101000111011001110111110011000010000110011001, 64'b0010011111101100111000010110110101111011100011100111101000110111,
          64'b0001010001000100010001110101000001110111011101100110100001101101, 64'b0000101000101100001101010000110000111001011000100110101110110011,
          64'b0000010100010111010111111000010101100100000100011000100111100001, 64'b0000001010001011110110000111100101110000101000001001100010100110,
          64'b0000000101000101111100010101010001000111010100010000101010111010, 64'b0000000010100010111110010100110100011011010000110000110011011011,
          64'b0000000001010001011111001011101011101100110000101010110011011110, 64'b0000000000101000101111100110000000000010010001101110100111101101,
          64'b0000000000010100010111110011000001010010101000000011001011011100, 64'b0000000000001010001011111001100000110011011111111011000110000110,
          64'b0000000000000101000101111100110000011011000001011100101111001001, 64'b0000000000000010100010111110011000001101101010111010010001000101,
          64'b0000000000000001010001011111001100000110110110101110100111101110, 64'b0000000000000000101000101111100110000011011011100001011111110000,
          64'b0000000000000000010100010111110011000001101101110010000001010111, 64'b0000000000000000001010001011111001100000110110111001001010110111,
          64'b0000000000000000000101000101111100110000011011011100100110101101, 64'b0000000000000000000010100010111110011000001101101110010011100000,
          64'b0000000000000000000001010001011111001100000110110111001001110001, 64'b0000000000000000000000101000101111100110000011011011100100111001,
          64'b0000000000000000000000010100010111110011000001101101110010011100, 64'b0000000000000000000000001010001011111001100000110110111001001110,
          64'b0000000000000000000000000101000101111100110000011011011100100111, 64'b0000000000000000000000000010100010111110011000001101101110010011,
          64'b0000000000000000000000000001010001011111001100000110110111001001, 64'b0000000000000000000000000000101000101111100110000011011011100100,
          64'b0000000000000000000000000000010100010111110011000001101101110010, 64'b0000000000000000000000000000001010001011111001100000110110111001,
          64'b0000000000000000000000000000000101000101111100110000011011011100, 64'b0000000000000000000000000000000010100010111110011000001101101110,
          64'b0000000000000000000000000000000001010001011111001100000110110111, 64'b0000000000000000000000000000000000101000101111100110000011011011,
          64'b0000000000000000000000000000000000010100010111110011000001101101, 64'b0000000000000000000000000000000000001010001011111001100000110110,
          64'b0000000000000000000000000000000000000101000101111100110000011011, 64'b0000000000000000000000000000000000000010100010111110011000001101,
          64'b0000000000000000000000000000000000000001010001011111001100000110, 64'b0000000000000000000000000000000000000000101000101111100110000011,
          64'b0000000000000000000000000000000000000000010100010111110011000001, 64'b0000000000000000000000000000000000000000001010001011111001100000,
          64'b0000000000000000000000000000000000000000000101000101111100110000, 64'b0000000000000000000000000000000000000000000010100010111110011000,
          64'b0000000000000000000000000000000000000000000001010001011111001100, 64'b0000000000000000000000000000000000000000000000101000101111100110,
          64'b0000000000000000000000000000000000000000000000010100010111110011, 64'b0000000000000000000000000000000000000000000000001010001011111001,
          64'b0000000000000000000000000000000000000000000000000101000101111100, 64'b0000000000000000000000000000000000000000000000000010100010111110,
          64'b0000000000000000000000000000000000000000000000000001010001011111, 64'b0000000000000000000000000000000000000000000000000000101000101111,
          64'b0000000000000000000000000000000000000000000000000000010100010111, 64'b0000000000000000000000000000000000000000000000000000001010001011,
          64'b0000000000000000000000000000000000000000000000000000000101000101, 64'b0000000000000000000000000000000000000000000000000000000010100010,
          64'b0000000000000000000000000000000000000000000000000000000001010001, 64'b0000000000000000000000000000000000000000000000000000000000101000,
          64'b0000000000000000000000000000000000000000000000000000000000010100, 64'b0000000000000000000000000000000000000000000000000000000000001010,
          64'b0000000000000000000000000000000000000000000000000000000000000101, 64'b0000000000000000000000000000000000000000000000000000000000000010,
          64'b0000000000000000000000000000000000000000000000000000000000000001, 64'b0000000000000000000000000000000000000000000000000000000000000000,
          64'b0000000000000000000000000000000000000000000000000000000000000000, {reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg
          , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_2mi_sva
          <= z_out_20[42:0];
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_x_2mi_sva
          <= operator_43_4_true_AC_TRN_AC_WRAP_4_rshift_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_6_4
          <= 3'b000;
    end
    else if ( ((fsm_output[13]) | (fsm_output[11]) | (fsm_output[6]) | (fsm_output[12]))
        & scatter_wen ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_6_4
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_rgt[6:4];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0
          <= 4'b0000;
    end
    else if ( ((fsm_output[11]) | (fsm_output[6]) | (fsm_output[13])) & scatter_wen
        ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_mux_rgt[3:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_37
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_36
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_32_31
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_24
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_23
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_18_17
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_15_14
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_9
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_8
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_7
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_6
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_4_0
          <= 5'b00000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_29
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_32_31
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_18_17
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_15_14
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_4_0
          <= 5'b00000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_35
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_34
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_32
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_31
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_18
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_17
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_15
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_14
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_0
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_37
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_36
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_32_31
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_24
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_23
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_18_17
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_15_14
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_9
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_8
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_7
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_6
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_4_0
          <= 5'b00000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_29
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_28
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_27
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_22
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_21
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_20
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_0
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_32_31
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_4_0
          <= 5'b00000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_35
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_34
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_32
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_31
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_29_27
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_22_20
          <= 3'b000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_18
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_17
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_15
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_14
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_0
          <= 1'b0;
    end
    else if ( and_2512_cse ) begin
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0
          <= ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_rgt[3:0];
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1}),
          (z_out_12[42:39]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_38
          <= MUX_s_1_2_2(z_out_1_33, (z_out_12[38]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_37
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[37]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_36
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[36]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_35_34
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_12[35:34]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_33
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[33]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_32_31
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_12[32:31]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_30
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[30]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(({{2{z_out_1_33}}, z_out_1_33}), (z_out_12[29:27]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_26
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[26]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_25
          <= MUX_s_1_2_2(z_out_1_33, (z_out_12[25]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_24
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[24]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_23
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[23]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(({{2{z_out_1_33}}, z_out_1_33}), (z_out_12[22:20]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[19]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_18_17
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_12[18:17]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_16
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[16]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_15_14
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_12[15:14]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_13
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[13]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_12
          <= MUX_s_1_2_2(z_out_1_33, (z_out_12[12]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_11
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[11]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_10
          <= MUX_s_1_2_2(z_out_1_33, (z_out_12[10]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_9
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[9]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_8
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[8]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_7
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[7]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_6
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_12[6]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_5
          <= MUX_s_1_2_2(z_out_1_33, (z_out_12[5]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_4_0
          <= MUX_v_5_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0}),
          (z_out_12[4:0]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_38
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[38]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_29
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[29]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_5
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[5]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28}),
          (z_out_16[42:39]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_35_34
          <= MUX_v_2_2_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27}),
          (z_out_16[35:34]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_32_31
          <= MUX_v_2_2_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26}),
          (z_out_16[32:31]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(({{2{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25}),
          (z_out_16[29:27]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(({{2{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9}),
          (z_out_16[22:20]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_18_17
          <= MUX_v_2_2_2(({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8}),
          (z_out_16[18:17]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_15_14
          <= MUX_v_2_2_2(({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7}),
          (z_out_16[15:14]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_4_0
          <= MUX_v_5_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14}),
          (z_out_16[4:0]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_38
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[38]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_35
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[35]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_34
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[34]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_32
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[32]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_31
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[31]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1,
          (z_out_10[29:27]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_25
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[25]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1,
          (z_out_10[22:20]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_18
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[18]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_17
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[17]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_15
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[15]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_14
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[14]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_12
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[12]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_10
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[10]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_5
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[5]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_0
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_10[0]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42
          <= MUX1HOT_v_3_3_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0}),
          (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6[44:42]),
          (z_out_7[44:42]), {(fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1}),
          (z_out_11[42:39]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_38
          <= MUX_s_1_2_2(z_out_1_33, (z_out_11[38]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_37
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[37]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_36
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[36]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_35_34
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_11[35:34]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_33
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[33]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_32_31
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_11[32:31]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_30
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[30]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(({{2{z_out_1_33}}, z_out_1_33}), (z_out_11[29:27]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_26
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[26]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_25
          <= MUX_s_1_2_2(z_out_1_33, (z_out_11[25]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_24
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[24]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_23
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[23]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(({{2{z_out_1_33}}, z_out_1_33}), (z_out_11[22:20]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_19
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[19]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_18_17
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_11[18:17]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_16
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[16]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_15_14
          <= MUX_v_2_2_2(({{1{z_out_1_33}}, z_out_1_33}), (z_out_11[15:14]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_13
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[13]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_12
          <= MUX_s_1_2_2(z_out_1_33, (z_out_11[12]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_11
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[11]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_10
          <= MUX_s_1_2_2(z_out_1_33, (z_out_11[10]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_9
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[9]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_8
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[8]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_7
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[7]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_6
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19_1,
          (z_out_11[6]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_5
          <= MUX_s_1_2_2(z_out_1_33, (z_out_11[5]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_4_0
          <= MUX_v_5_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0}),
          (z_out_11[4:0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_or_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42
          <= MUX1HOT_v_3_3_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17}),
          (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6[44:42]),
          (z_out_8[44:42]), {(fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_38
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[38]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_29
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[29]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_28
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[28]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_27
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[27]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_25
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[25]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_22
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[22]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_21
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[21]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_20
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[20]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_12
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[12]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_10
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[10]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_5
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[5]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_0
          <= MUX_s_1_2_2(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_13[0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42
          <= MUX1HOT_v_3_3_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42}),
          (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6[44:42]),
          (z_out_6[44:42]), {(fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(({{3{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28}),
          (z_out_15[42:39]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_35_34
          <= MUX_v_2_2_2(({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24}),
          (z_out_15[35:34]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_32_31
          <= MUX_v_2_2_2(({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22}),
          (z_out_15[32:31]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(({{2{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20}),
          (z_out_15[29:27]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(({{2{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16}),
          (z_out_15[22:20]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_4_0
          <= MUX_v_5_2_2(({{3{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0}),
          (z_out_15[4:0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42
          <= MUX1HOT_v_3_3_2(({{1{ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0[1]}},
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0}),
          (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6[44:42]),
          (z_out_9[44:42]), {(fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt
          , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_38
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[38]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_35
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[35]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_34
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[34]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_32
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[32]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_31
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[31]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_29_27
          <= MUX_v_3_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1,
          (z_out_17[29:27]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_25
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[25]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_22_20
          <= MUX_v_3_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1,
          (z_out_17[22:20]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_18
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[18]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_17
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[17]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_15
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[15]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_14
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[14]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_12
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[12]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_10
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[10]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_5
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[5]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_0
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20_1[2]),
          (z_out_17[0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_19
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_38
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_5
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_37
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_36
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_9
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_6
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_8
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_7
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_10
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_33
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_11
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_12
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_30
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_13
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_26
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_16
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_24
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_23
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_32_31
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_15_14
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_18_17
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_35_34
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_32_31
          <= 2'b00;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_9_cse
        ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_19
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[19]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_38
          <= MUX_s_1_2_2(z_out_1_33, (z_out_16[38]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_5
          <= MUX_s_1_2_2(z_out_1_33, (z_out_16[5]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_37
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[37]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_36
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[36]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_9
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[9]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_6
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[6]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_8
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[8]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_7
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[7]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_10
          <= MUX_s_1_2_2(z_out_1_33, (z_out_16[10]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_33
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[33]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_11
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[11]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_12
          <= MUX_s_1_2_2(z_out_1_33, (z_out_16[12]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_30
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[30]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_13
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[13]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_26
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[26]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_16
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[16]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_25
          <= MUX_s_1_2_2(z_out_1_33, (z_out_16[25]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_24
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[24]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_23
          <= MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          (z_out_16[23]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_13[18:17]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_35_34
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_13[35:34]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_32_31
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_13[32:31]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_15_14
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_13[15:14]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_18_17
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_14[18:17]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_35_34
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_14[35:34]), fsm_output[13]);
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_32_31
          <= MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1,
          (z_out_14[32:31]), fsm_output[13]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_0
          <= 1'b0;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_29_cse
        ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse
          <= ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1[1];
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_0
          <= MUX_s_1_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17_1[1]),
          (z_out_4[28]), fsm_output[17]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0
          <= 2'b00;
    end
    else if ( and_2513_cse ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42
          <= MUX_v_2_2_2(2'b00, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_5_nl),
          (not_340_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0
          <= MUX_v_2_2_2(2'b00, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_4_nl),
          (not_339_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28
          <= 1'b0;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17
          <= 2'b00;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_and_6_cse
        ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25
          <= MUX1HOT_s_1_3_2(z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[25]), {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27
          <= MUX1HOT_s_1_3_2(z_out_1_33, reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[27]), {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28
          <= MUX1HOT_s_1_3_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
          reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_38_cse,
          (z_out_14[28]), {(fsm_output[9]) , (fsm_output[11]) , (fsm_output[13])});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14
          <= MUX1HOT_v_2_3_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0,
          ({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12}),
          (z_out_15[15:14]), {(fsm_output[9]) , (fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17
          <= MUX1HOT_v_2_3_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0,
          ({{1{ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14}},
          ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14}),
          (z_out_15[18:17]), {(fsm_output[9]) , (fsm_output[11]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21 <= 12'b000000000000;
    end
    else if ( ((fsm_output[15]) | (fsm_output[16]) | (fsm_output[17]) | (fsm_output[18])
        | (fsm_output[14]) | (fsm_output[10])) & scatter_wen ) begin
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21 <= lambertianScatter_rand_unit_run_phi_mux1h_2_rgt[32:21];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0 <= 21'b000000000000000000000;
    end
    else if ( ((fsm_output[14]) | (fsm_output[10])) & scatter_wen ) begin
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0 <= lambertianScatter_rand_unit_run_phi_mux1h_2_rgt[20:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_9_6
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_37_36
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_24_23
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_9_6
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_4_1
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0
          <= 42'b000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_37_36
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_24_23
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_9_6
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_4_1
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0
          <= 42'b000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_42_39
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_37_36
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_24_23
          <= 2'b00;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_9_6
          <= 4'b0000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_4_1
          <= 4'b0000;
    end
    else if ( and_2517_cse ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_9_6
          <= MUX_v_4_2_2(4'b0000, (z_out_14[9:6]), (not_335_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(4'b0000, (z_out_10[42:39]), (not_334_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_37_36
          <= MUX_v_2_2_2(2'b00, (z_out_10[37:36]), (not_333_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_24_23
          <= MUX_v_2_2_2(2'b00, (z_out_10[24:23]), (not_329_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_9_6
          <= MUX_v_4_2_2(4'b0000, (z_out_10[9:6]), (not_324_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_4_1
          <= MUX_v_4_2_2(4'b0000, (z_out_10[4:1]), (not_323_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0
          <= MUX_v_42_2_2(42'b000000000000000000000000000000000000000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_1_nl),
          (not_321_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(4'b0000, (z_out_13[42:39]), (not_318_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_37_36
          <= MUX_v_2_2_2(2'b00, (z_out_13[37:36]), (not_317_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_24_23
          <= MUX_v_2_2_2(2'b00, (z_out_13[24:23]), (not_313_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_9_6
          <= MUX_v_4_2_2(4'b0000, (z_out_13[9:6]), (not_308_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_4_1
          <= MUX_v_4_2_2(4'b0000, (z_out_13[4:1]), (not_307_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0
          <= MUX_v_42_2_2(42'b000000000000000000000000000000000000000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_nl),
          (not_304_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_42_39
          <= MUX_v_4_2_2(4'b0000, (z_out_17[42:39]), (not_303_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_37_36
          <= MUX_v_2_2_2(2'b00, (z_out_17[37:36]), (not_302_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_24_23
          <= MUX_v_2_2_2(2'b00, (z_out_17[24:23]), (not_298_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_9_6
          <= MUX_v_4_2_2(4'b0000, (z_out_17[9:6]), (not_293_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_4_1
          <= MUX_v_4_2_2(4'b0000, (z_out_17[4:1]), (not_292_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva
          <= 6'b000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva
          <= 6'b000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva
          <= 6'b000000;
    end
    else if ( and_2523_cse ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva
          <= MUX_v_6_2_2(6'b000000, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva_3,
          (not_322_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva
          <= MUX_v_6_2_2(6'b000000, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva_2,
          (not_320_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva
          <= MUX_v_6_2_2(6'b000000, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva_2,
          (not_305_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36
          <= 6'b000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36
          <= 6'b000000;
    end
    else if ( and_2527_cse ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36
          <= MUX_v_6_2_2(6'b000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_1_nl),
          (not_533_nl));
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36
          <= MUX_v_6_2_2(6'b000000, (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_nl),
          (not_534_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_y_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
    end
    else if ( scatter_wen & and_dcpl_5 & and_8_cse ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_y_2mi_sva
          <= operator_43_4_true_AC_TRN_AC_WRAP_7_rshift_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs
          <= 1'b0;
    end
    else if ( scatter_wen & ((fsm_output[12]) | or_tmp_78 | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs_mx0c2)
        ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs
          <= MUX1HOT_s_1_3_2((z_out_7[45]), (else_else_and_1_nl), (ray_in_crt_sva[165]),
          {(fsm_output[12]) , or_tmp_78 , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs_mx0c2});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_atan_pi_2mi_return_69_28_sva <= 42'b000000000000000000000000000000000000000000;
      ac_math_atan_pi_2mi_return_1_69_28_sva <= 42'b000000000000000000000000000000000000000000;
      ac_math_atan_pi_2mi_return_2_69_28_sva <= 42'b000000000000000000000000000000000000000000;
      ac_math_atan_pi_2mi_return_3_69_28_sva <= 42'b000000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_d_a_and_cse
        ) begin
      ac_math_atan_pi_2mi_return_69_28_sva <= MUX_v_42_37_2(42'b100000000000000000000000000000000000000000,
          42'b010010111001000000010100011101100111011111, 42'b001001111110110011100001011011010111101110,
          42'b000101000100010001000111010100000111011101, 42'b000010100010110000110101000011000011100101,
          42'b000001010001011101011111100001010110010000, 42'b000000101000101111011000011110010111000010,
          42'b000000010100010111110001010101000100011101, 42'b000000001010001011111001010011010001101101,
          42'b000000000101000101111100101110101110110011, 42'b000000000010100010111110011000000000001001,
          42'b000000000001010001011111001100000101001010, 42'b000000000000101000101111100110000011001101,
          42'b000000000000010100010111110011000001101100, 42'b000000000000001010001011111001100000110110,
          42'b000000000000000101000101111100110000011011, 42'b000000000000000010100010111110011000001101,
          42'b000000000000000001010001011111001100000110, 42'b000000000000000000101000101111100110000011,
          42'b000000000000000000010100010111110011000001, 42'b000000000000000000001010001011111001100000,
          42'b000000000000000000000101000101111100110000, 42'b000000000000000000000010100010111110011000,
          42'b000000000000000000000001010001011111001100, 42'b000000000000000000000000101000101111100110,
          42'b000000000000000000000000010100010111110011, 42'b000000000000000000000000001010001011111001,
          42'b000000000000000000000000000101000101111100, 42'b000000000000000000000000000010100010111110,
          42'b000000000000000000000000000001010001011111, 42'b000000000000000000000000000000101000101111,
          42'b000000000000000000000000000000010100010111, 42'b000000000000000000000000000000001010001011,
          42'b000000000000000000000000000000000101000101, 42'b000000000000000000000000000000000010100010,
          42'b000000000000000000000000000000000001010001, 42'b000000000000000000000000000000000000101000,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_5_0_sva);
      ac_math_atan_pi_2mi_return_1_69_28_sva <= MUX_v_42_37_2(42'b100000000000000000000000000000000000000000,
          42'b010010111001000000010100011101100111011111, 42'b001001111110110011100001011011010111101110,
          42'b000101000100010001000111010100000111011101, 42'b000010100010110000110101000011000011100101,
          42'b000001010001011101011111100001010110010000, 42'b000000101000101111011000011110010111000010,
          42'b000000010100010111110001010101000100011101, 42'b000000001010001011111001010011010001101101,
          42'b000000000101000101111100101110101110110011, 42'b000000000010100010111110011000000000001001,
          42'b000000000001010001011111001100000101001010, 42'b000000000000101000101111100110000011001101,
          42'b000000000000010100010111110011000001101100, 42'b000000000000001010001011111001100000110110,
          42'b000000000000000101000101111100110000011011, 42'b000000000000000010100010111110011000001101,
          42'b000000000000000001010001011111001100000110, 42'b000000000000000000101000101111100110000011,
          42'b000000000000000000010100010111110011000001, 42'b000000000000000000001010001011111001100000,
          42'b000000000000000000000101000101111100110000, 42'b000000000000000000000010100010111110011000,
          42'b000000000000000000000001010001011111001100, 42'b000000000000000000000000101000101111100110,
          42'b000000000000000000000000010100010111110011, 42'b000000000000000000000000001010001011111001,
          42'b000000000000000000000000000101000101111100, 42'b000000000000000000000000000010100010111110,
          42'b000000000000000000000000000001010001011111, 42'b000000000000000000000000000000101000101111,
          42'b000000000000000000000000000000010100010111, 42'b000000000000000000000000000000001010001011,
          42'b000000000000000000000000000000000101000101, 42'b000000000000000000000000000000000010100010,
          42'b000000000000000000000000000000000001010001, 42'b000000000000000000000000000000000000101000,
          reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg);
      ac_math_atan_pi_2mi_return_2_69_28_sva <= MUX_v_42_37_2(42'b100000000000000000000000000000000000000000,
          42'b010010111001000000010100011101100111011111, 42'b001001111110110011100001011011010111101110,
          42'b000101000100010001000111010100000111011101, 42'b000010100010110000110101000011000011100101,
          42'b000001010001011101011111100001010110010000, 42'b000000101000101111011000011110010111000010,
          42'b000000010100010111110001010101000100011101, 42'b000000001010001011111001010011010001101101,
          42'b000000000101000101111100101110101110110011, 42'b000000000010100010111110011000000000001001,
          42'b000000000001010001011111001100000101001010, 42'b000000000000101000101111100110000011001101,
          42'b000000000000010100010111110011000001101100, 42'b000000000000001010001011111001100000110110,
          42'b000000000000000101000101111100110000011011, 42'b000000000000000010100010111110011000001101,
          42'b000000000000000001010001011111001100000110, 42'b000000000000000000101000101111100110000011,
          42'b000000000000000000010100010111110011000001, 42'b000000000000000000001010001011111001100000,
          42'b000000000000000000000101000101111100110000, 42'b000000000000000000000010100010111110011000,
          42'b000000000000000000000001010001011111001100, 42'b000000000000000000000000101000101111100110,
          42'b000000000000000000000000010100010111110011, 42'b000000000000000000000000001010001011111001,
          42'b000000000000000000000000000101000101111100, 42'b000000000000000000000000000010100010111110,
          42'b000000000000000000000000000001010001011111, 42'b000000000000000000000000000000101000101111,
          42'b000000000000000000000000000000010100010111, 42'b000000000000000000000000000000001010001011,
          42'b000000000000000000000000000000000101000101, 42'b000000000000000000000000000000000010100010,
          42'b000000000000000000000000000000000001010001, 42'b000000000000000000000000000000000000101000,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_i_5_0_sva);
      ac_math_atan_pi_2mi_return_3_69_28_sva <= MUX_v_42_37_2(42'b100000000000000000000000000000000000000000,
          42'b010010111001000000010100011101100111011111, 42'b001001111110110011100001011011010111101110,
          42'b000101000100010001000111010100000111011101, 42'b000010100010110000110101000011000011100101,
          42'b000001010001011101011111100001010110010000, 42'b000000101000101111011000011110010111000010,
          42'b000000010100010111110001010101000100011101, 42'b000000001010001011111001010011010001101101,
          42'b000000000101000101111100101110101110110011, 42'b000000000010100010111110011000000000001001,
          42'b000000000001010001011111001100000101001010, 42'b000000000000101000101111100110000011001101,
          42'b000000000000010100010111110011000001101100, 42'b000000000000001010001011111001100000110110,
          42'b000000000000000101000101111100110000011011, 42'b000000000000000010100010111110011000001101,
          42'b000000000000000001010001011111001100000110, 42'b000000000000000000101000101111100110000011,
          42'b000000000000000000010100010111110011000001, 42'b000000000000000000001010001011111001100000,
          42'b000000000000000000000101000101111100110000, 42'b000000000000000000000010100010111110011000,
          42'b000000000000000000000001010001011111001100, 42'b000000000000000000000000101000101111100110,
          42'b000000000000000000000000010100010111110011, 42'b000000000000000000000000001010001011111001,
          42'b000000000000000000000000000101000101111100, 42'b000000000000000000000000000010100010111110,
          42'b000000000000000000000000000001010001011111, 42'b000000000000000000000000000000101000101111,
          42'b000000000000000000000000000000010100010111, 42'b000000000000000000000000000000001010001011,
          42'b000000000000000000000000000000000101000101, 42'b000000000000000000000000000000000010100010,
          42'b000000000000000000000000000000000001010001, 42'b000000000000000000000000000000000000101000,
          ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_i_5_0_sva);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_y_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
    end
    else if ( ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_and_cse
        ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_sva
          <= operator_43_4_true_AC_TRN_AC_WRAP_1_rshift_itm;
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_y_2mi_sva
          <= operator_43_4_true_AC_TRN_AC_WRAP_5_rshift_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_x_2mi_sva
          <= 43'b0000000000000000000000000000000000000000000;
    end
    else if ( scatter_wen & and_dcpl_5 & and_dcpl_18 & (~ else_unequal_tmp) ) begin
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_x_2mi_sva
          <= operator_43_4_true_AC_TRN_AC_WRAP_6_rshift_itm;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mux_21_itm <= 21'b000000000000000000000;
    end
    else if ( scatter_wen & (or_tmp_111 | and_352_cse) ) begin
      mux_21_itm <= MUX_v_21_2_2((hit_in_crt_sva_171_0[62:42]), (ray_in_crt_sva[62:42]),
          and_352_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_lambertianScatter_add_run_acc_psp_ftd <= 26'b00000000000000000000000000;
    end
    else if ( scatter_wen & (~ or_dcpl_30) & (fsm_output[16]) ) begin
      reg_lambertianScatter_add_run_acc_psp_ftd <= z_out_18[26:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_lambertianScatter_add_run_acc_3_psp_ftd <= 26'b00000000000000000000000000;
    end
    else if ( scatter_wen & (~ or_dcpl_30) & (fsm_output[17]) ) begin
      reg_lambertianScatter_add_run_acc_3_psp_ftd <= z_out_18[26:1];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2
          <= 8'b00000000;
    end
    else if ( scatter_wen & (~((fsm_output[17]) | (fsm_output[15]) | or_dcpl_73))
        ) begin
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2
          <= MUX_v_8_2_2((operator_43_4_true_AC_TRN_AC_WRAP_2_rshift_itm[14:7]),
          (z_out_10[14:7]), fsm_output[13]);
    end
  end
  assign lambertianScatter_run_mux_nl = MUX_v_26_2_2(reg_lambertianScatter_add_run_acc_psp_ftd,
      (signext_26_25(hit_in_crt_sva_171_0[88:64])), lambertianScatter_run_land_1_lpi_1_dfm_mx2);
  assign lambertianScatter_run_mux_1_nl = MUX_v_26_2_2(reg_lambertianScatter_add_run_acc_3_psp_ftd,
      (signext_26_25(hit_in_crt_sva_171_0[114:90])), lambertianScatter_run_land_1_lpi_1_dfm_mx2);
  assign lambertianScatter_run_mux_2_nl = MUX_v_26_2_2((lambertianScatter_add_run_acc_4_psp_sva[26:1]),
      (signext_26_25(hit_in_crt_sva_171_0[140:116])), lambertianScatter_run_land_1_lpi_1_dfm_mx2);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_4_nl
      = MUX1HOT_s_1_5_2((z_out_3[28]), rand_unit_random2_run_x3_28_sva_mx0w0, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19_mx1w2,
      (z_out_14[19]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
      , or_tmp_208 , (fsm_output[9]) , (fsm_output[13])});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_8_nl
      = MUX1HOT_s_1_5_2((z_out_3[24]), rand_unit_random2_run_x3_24_sva_mx0w0, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24,
      z_out_1_33, (z_out_14[16]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
      , or_tmp_208 , (fsm_output[9]) , (fsm_output[13])});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_17_nl
      = MUX1HOT_s_1_5_2((z_out_3[22]), rand_unit_random2_run_x3_22_sva_mx0w0, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22,
      z_out_1_33, (z_out_14[13]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
      , or_tmp_208 , (fsm_output[9]) , (fsm_output[13])});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux1h_41_nl
      = MUX1HOT_s_1_5_2((z_out_3[16]), rand_unit_random2_run_x3_16_sva_mx0w0, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16,
      z_out_1_33, (z_out_14[11]), {ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_43_cse
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_and_44_cse
      , or_tmp_208 , (fsm_output[9]) , (fsm_output[13])});
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm
      + z_out_20 + 69'b000000000000000000000000000000000000000000000000000000000000000000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux1h_89_nl
      = MUX1HOT_s_1_3_2(z_out_1_33, ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26,
      (z_out_14[26]), {(fsm_output[9]) , or_tmp_516 , (fsm_output[13])});
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_33_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33,
      (z_out_14[33]), fsm_output[13]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_32_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30,
      (z_out_14[30]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33,
      (z_out_10[33]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30,
      (z_out_10[30]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_7_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26,
      (z_out_10[26]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19,
      (z_out_10[19]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16,
      (z_out_10[16]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13,
      (z_out_10[13]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_2_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11,
      (z_out_10[11]), fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_or_3_nl
      = (fsm_output[12]) | (fsm_output[14]);
  assign and_202_nl = (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm)
      & ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_16_nl
      = MUX1HOT_v_36_4_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0,
      (z_out_8[35:0]), (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6[35:0]),
      (z_out_16[42:7]), {(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_or_3_nl)
      , (and_202_nl) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_4_ssc
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_11_cse});
  assign not_319_nl = ~ (fsm_output[11]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_6_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33,
      (z_out_13[33]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_5_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30,
      (z_out_13[30]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_4_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26,
      (z_out_13[26]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_3_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19,
      (z_out_13[19]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_2_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16,
      (z_out_13[16]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_1_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13,
      (z_out_13[13]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11,
      (z_out_13[11]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_or_3_rgt);
  assign and_204_nl = (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_and_itm)
      & ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1
      & (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux1h_15_nl
      = MUX1HOT_v_36_5_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0,
      (z_out_6[35:0]), (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6[35:0]),
      (z_out_14[42:7]), (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva[42:7]),
      {(fsm_output[12]) , (and_204_nl) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_1_ssc
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_11_cse
      , (fsm_output[14])});
  assign not_306_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_10_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33,
      (z_out_17[33]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_9_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30,
      (z_out_17[30]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_8_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26,
      (z_out_17[26]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_6_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19,
      (z_out_17[19]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_5_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16,
      (z_out_17[16]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_4_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13,
      (z_out_17[13]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_mux_3_nl
      = MUX_s_1_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11,
      (z_out_17[11]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_or_12_cse);
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl
      = conv_u2s_6_7(z_out_3[6:1]) + 7'b1011111;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_nl[6:0];
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva
      + z_out_20 + 69'b000000000000000000000000000000000000000000000000000000000000000000001;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_1_nl[68:0];
  assign nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva +
      z_out_20;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl
      = nl_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_3_nl[68:0];
  assign not_341_nl = ~ (fsm_output[5]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_or_nl
      = ((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm[68])
      & (z_out_5[69])) | (~((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_mux_2_itm[68])
      | (z_out_5[69])));
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_2_nor_nl
      = ~((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_lpi_1_dfm_64_0_mx0[31:0]!=32'b00000000000000000000000000000000));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_5_nl
      = MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0,
      (z_out_14[37:36]), fsm_output[13]);
  assign not_340_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_4_nl
      = MUX_v_2_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42_mx1w0,
      (z_out_14[24:23]), fsm_output[13]);
  assign not_339_nl = ~ (fsm_output[11]);
  assign not_335_nl = ~ (fsm_output[11]);
  assign not_334_nl = ~ (fsm_output[11]);
  assign not_333_nl = ~ (fsm_output[11]);
  assign not_329_nl = ~ (fsm_output[11]);
  assign not_324_nl = ~ (fsm_output[11]);
  assign not_323_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_1_nl
      = MUX_v_42_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_sva_6[41:0]),
      (z_out_7[41:0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt);
  assign not_321_nl = ~ (fsm_output[11]);
  assign not_318_nl = ~ (fsm_output[11]);
  assign not_317_nl = ~ (fsm_output[11]);
  assign not_313_nl = ~ (fsm_output[11]);
  assign not_308_nl = ~ (fsm_output[11]);
  assign not_307_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_mux_nl
      = MUX_v_42_2_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_sva_6[41:0]),
      (z_out_9[41:0]), ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt);
  assign not_304_nl = ~ (fsm_output[11]);
  assign not_303_nl = ~ (fsm_output[11]);
  assign not_302_nl = ~ (fsm_output[11]);
  assign not_298_nl = ~ (fsm_output[11]);
  assign not_293_nl = ~ (fsm_output[11]);
  assign not_292_nl = ~ (fsm_output[11]);
  assign not_322_nl = ~ (fsm_output[11]);
  assign not_320_nl = ~ (fsm_output[11]);
  assign not_305_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_1_nl
      = MUX_v_6_2_2((z_out_8[41:36]), (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_sva_6[41:36]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_4_ssc);
  assign not_533_nl = ~ (fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_mux_nl
      = MUX_v_6_2_2((z_out_6[41:36]), (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_sva_6[41:36]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_and_1_ssc);
  assign not_534_nl = ~ (fsm_output[11]);
  assign else_else_and_1_nl = (ray_in_crt_sva[165]) & else_unequal_tmp;
  assign else_else_mux1h_1_nl = MUX1HOT_v_27_3_2((accumalated_color_chan_in_crt_sva[53:27]),
      (accumalated_color_chan_in_crt_sva[80:54]), (accumalated_color_chan_in_crt_sva[26:0]),
      {(fsm_output[4]) , (fsm_output[3]) , (fsm_output[5])});
  assign nl_z_out = else_if_mul_cmp_z_oreg + (else_else_mux1h_1_nl);
  assign z_out = nl_z_out[26:0];
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_32_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_31), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[11])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_33_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_30), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[10])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_34_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_29), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[9])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_35_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_28), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[8])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_36_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_27), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[7])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_37_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_26), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[6])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_38_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_25), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[5])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_39_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_24), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[4])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_40_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_23), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[3])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_41_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_22), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[2])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_42_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_21), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[1])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_43_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_20), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[0])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_44_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_19), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[20])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_45_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_18), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[19])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_46_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_17), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[18])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_47_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_16), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[17])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_48_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_15), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[16])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_49_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_14), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[15])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_50_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_13), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[14])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_51_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_12), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[13])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_52_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_11), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[12])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_53_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_10), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[11])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_54_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_9), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[10])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_55_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_8), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[9])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_56_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_7), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[8])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_57_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_6), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[7])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_58_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x3_sva_5), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[6])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_59_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x2_12_0_sva_4), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[5])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_60_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x2_12_0_sva_3), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[4])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_61_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x2_12_0_sva_2), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[3])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_62_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x2_12_0_sva_1), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[2])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_63_nl
      = MUX_s_1_2_2((~ rand_unit_random1_run_x2_12_0_sva_0), (~ (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[1])),
      fsm_output[11]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_nand_1_nl
      = ~((lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0[0]) & (fsm_output[11]));
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl
      = conv_s2u_33_34({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_32_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_33_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_34_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_35_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_36_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_37_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_38_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_39_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_40_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_41_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_42_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_43_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_44_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_45_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_46_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_47_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_48_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_49_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_50_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_51_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_52_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_53_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_54_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_55_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_56_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_57_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_58_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_59_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_60_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_61_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_62_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_mux_63_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_nand_1_nl)})
      + 34'b0010000000000000000000000000000001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl[33:0];
  assign z_out_1_33 = readslicef_34_1_33((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_if_acc_nl));
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_31_nl
      = ~(lambertianScatter_state2_17_sva ^ xor_cse_9);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_31_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_31_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_32_nl
      = MUX_s_1_2_2((~ xor_cse_11), reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_32_nl
      = ~(lambertianScatter_state2_10_sva ^ xor_cse_3);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_33_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_32_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_33_nl
      = ~(lambertianScatter_state2_14_sva ^ xor_cse_14);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_34_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_33_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_34_nl
      = ~(lambertianScatter_state2_13_sva ^ xor_cse_17);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_35_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_34_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_35_nl
      = ~(lambertianScatter_state2_12_sva ^ xor_cse_18);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_36_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_35_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_36_nl
      = ~(lambertianScatter_state2_24_sva ^ lambertianScatter_state2_11_sva ^ lambertianScatter_state2_19_sva
      ^ lambertianScatter_state2_6_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_37_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_36_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_37_nl
      = ~(lambertianScatter_state2_23_sva ^ lambertianScatter_state2_10_sva ^ lambertianScatter_state2_18_sva
      ^ lambertianScatter_state2_5_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_38_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_37_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_38_nl
      = ~(lambertianScatter_state2_22_sva ^ lambertianScatter_state2_9_sva ^ lambertianScatter_state2_17_sva
      ^ lambertianScatter_state2_4_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_39_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_38_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_39_nl
      = ~(lambertianScatter_state2_21_sva ^ lambertianScatter_state2_8_sva ^ lambertianScatter_state2_16_sva
      ^ lambertianScatter_state2_3_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_40_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_39_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_40_nl
      = ~(lambertianScatter_state2_20_sva ^ lambertianScatter_state2_7_sva ^ lambertianScatter_state2_15_sva
      ^ lambertianScatter_state2_2_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_41_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_40_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_41_nl
      = ~(lambertianScatter_state2_6_sva ^ lambertianScatter_state2_14_sva ^ xor_cse_20);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_42_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_41_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_42_nl
      = ~(lambertianScatter_state2_18_sva ^ lambertianScatter_state2_5_sva ^ xor_cse_15);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_43_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_42_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_43_nl
      = ~(lambertianScatter_state2_16_sva ^ xor_cse_2);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_44_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_43_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_44_nl
      = ~(lambertianScatter_state2_11_sva ^ xor_cse_19);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_45_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_44_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_45_nl
      = ~(lambertianScatter_state2_10_sva ^ xor_cse_10);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_46_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_45_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_46_nl
      = ~(xor_cse_12 ^ xor_cse_13);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_47_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_46_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_47_nl
      = ~(xor_cse_15 ^ xor_cse_16);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_48_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_47_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_48_nl
      = ~(lambertianScatter_state2_12_sva ^ lambertianScatter_state2_7_sva ^ xor_cse_11);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_49_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_48_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_49_nl
      = ~(lambertianScatter_state2_28_sva ^ lambertianScatter_state2_15_sva ^ xor_cse);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_50_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_49_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_50_nl
      = ~(lambertianScatter_state2_27_sva ^ lambertianScatter_state2_14_sva ^ xor_cse_1);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_51_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_50_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_51_nl
      = ~(lambertianScatter_state2_13_sva ^ lambertianScatter_state2_4_sva ^ xor_cse_4);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_52_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_51_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_52_nl
      = ~(lambertianScatter_state2_3_sva ^ lambertianScatter_state2_20_sva ^ xor_cse_6);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_53_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_52_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_53_nl
      = ~(lambertianScatter_state2_19_sva ^ lambertianScatter_state2_6_sva ^ xor_cse_8);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_54_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_53_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_54_nl
      = ~(lambertianScatter_state2_10_sva ^ lambertianScatter_state2_5_sva ^ xor_cse_7);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_55_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_54_nl),
      reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg,
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_55_nl
      = ~(lambertianScatter_state2_0_sva ^ lambertianScatter_state2_17_sva ^ xor_cse_5);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_56_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_55_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[5]),
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_56_nl
      = ~(lambertianScatter_state2_4_sva ^ lambertianScatter_state2_21_sva ^ lambertianScatter_state2_8_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_57_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_56_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[4]),
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_57_nl
      = ~(lambertianScatter_state2_3_sva ^ lambertianScatter_state2_20_sva ^ lambertianScatter_state2_7_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_58_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_57_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[3]),
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_58_nl
      = ~(lambertianScatter_state2_2_sva ^ lambertianScatter_state2_19_sva ^ lambertianScatter_state2_6_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_59_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_58_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[2]),
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_59_nl
      = ~(lambertianScatter_state2_1_sva ^ lambertianScatter_state2_18_sva ^ lambertianScatter_state2_5_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_60_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_59_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[1]),
      fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_60_nl
      = ~(lambertianScatter_state2_0_sva ^ lambertianScatter_state2_17_sva ^ lambertianScatter_state2_4_sva);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_61_nl
      = MUX_s_1_2_2((ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_xnor_60_nl),
      (reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg[0]),
      fsm_output[6]);
  assign nl_z_out_3 = conv_u2u_31_32({(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_31_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_32_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_33_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_34_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_35_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_36_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_37_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_38_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_39_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_40_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_41_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_42_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_43_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_44_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_45_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_46_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_47_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_48_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_49_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_50_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_51_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_52_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_53_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_54_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_55_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_56_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_57_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_58_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_59_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_60_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_if_mux_61_nl)})
      + 32'b00000000000000000000000000000001;
  assign z_out_3 = nl_z_out_3[31:0];
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_2_nl
      = lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_27 &
      or_1202_ssc;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_3_nl
      = MUX_v_20_2_2(20'b00000000000000000000, (lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0[26:7]),
      or_1202_ssc);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_2_nl
      = MUX_v_7_2_2(({reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_reg
      , reg_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_2_reg}),
      (lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0[6:0]),
      or_1202_ssc);
  assign nl_z_out_4 = conv_u2u_28_29({(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_2_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_and_3_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_mux_2_nl)})
      + 29'b11111111111111111111111111111;
  assign z_out_4 = nl_z_out_4[28:0];
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_4_nl
      = ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse
      | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_1_nl
      = MUX_v_69_2_2(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_1_sva,
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_sva, ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_4_nl);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_5_nl
      = (~(or_tmp_1118 | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse))
      | or_tmp_1119 | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse
      | (fsm_output[6]);
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_6_nl
      = or_tmp_1118 | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_2_cse;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_7_nl
      = or_tmp_1119 | ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_theta_and_1_cse;
  assign ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux1h_1_nl
      = MUX1HOT_v_69_3_2(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_sva,
      (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_sva),
      (~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_tn_sva),
      {(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_6_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_7_nl)
      , (fsm_output[6])});
  assign nl_acc_5_nl = conv_s2u_70_71({(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_1_nl)
      , (ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_5_nl)})
      + conv_s2u_70_71({(ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux1h_1_nl)
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[70:0];
  assign z_out_5 = readslicef_71_70_1((acc_5_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_33_nl
      = MUX_v_3_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_44_42,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_34_nl
      = MUX_v_6_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_41_36,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_35_nl
      = MUX_v_36_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_acc_a_lpi_1_dfm_1_35_0,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_36_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_29, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[41])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_37_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_28, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[40])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_38_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_27, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[39])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_39_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_26, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[38])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_40_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_25, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[37])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_41_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_24, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[36])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_42_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_23, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[35])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_43_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_22, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[34])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_44_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_21, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[33])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_45_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_20, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[32])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_46_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_19, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[31])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_47_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_18, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[30])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_48_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_17, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[29])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_49_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_16, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[28])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_50_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_15, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[27])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_51_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_14, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[26])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_52_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_13, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[25])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_53_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_12, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[24])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_54_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_11, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[23])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_55_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_10, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[22])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_56_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_9, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[21])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_57_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_8, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[20])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_58_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_7, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[19])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_59_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_6, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[18])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_60_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_5, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[17])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_61_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_4, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[16])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_62_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_3, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[15])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_63_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_2, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[14])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_64_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_1, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[13])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_65_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_0, (~ (ac_math_atan_pi_2mi_return_1_69_28_sva[12])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_not_61_nl
      = ~ (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_n000000
      = ~(MUX_v_12_2_2((ac_math_atan_pi_2mi_return_1_69_28_sva[11:0]), 12'b111111111111,
      (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_not_61_nl)));
  assign nl_acc_6_nl = conv_s2u_46_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_33_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_34_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_35_nl)
      , 1'b1}) + conv_s2u_45_47({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_1_cse
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_36_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_37_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_38_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_39_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_40_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_41_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_42_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_43_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_44_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_45_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_46_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_47_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_48_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_49_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_50_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_51_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_52_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_53_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_54_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_55_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_56_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_57_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_58_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_59_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_60_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_61_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_62_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_63_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_64_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_mux_65_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_n000000)
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[46:0];
  assign z_out_6 = readslicef_47_46_1((acc_6_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_32_nl
      = MUX_v_3_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_44_42,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_33_nl
      = MUX_v_42_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_lpi_1_dfm_1_41_0,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_34_nl
      = MUX_v_44_2_2(({lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21 ,
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0 , 11'b00000000000}),
      ({2'b11 , (~ ac_math_atan_pi_2mi_return_3_69_28_sva)}), fsm_output[13]);
  assign nl_acc_7_nl = conv_s2u_46_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_32_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_33_nl)
      , 1'b1}) + conv_s2u_45_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_34_nl)
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[46:0];
  assign z_out_7 = readslicef_47_46_1((acc_7_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_63_nl
      = MUX_v_3_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_44_42,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_64_nl
      = MUX_v_6_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_41_36,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_65_nl
      = MUX_v_36_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_acc_a_lpi_1_dfm_1_35_0,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_66_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_29, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[41])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_67_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_28, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[40])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_68_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_27, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[39])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_69_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_26, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[38])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_70_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_25, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[37])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_71_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_24, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[36])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_72_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_23, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[35])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_73_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_22, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[34])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_74_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_21, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[33])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_75_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_20, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[32])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_76_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_19, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[31])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_77_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_18, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[30])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_78_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_17, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[29])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_79_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_16, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[28])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_80_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_15, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[27])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_81_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_14, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[26])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_82_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_13, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[25])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_83_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_12, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[24])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_84_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_11, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[23])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_85_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_10, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[22])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_86_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_9, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[21])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_87_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_8, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[20])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_88_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_7, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[19])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_89_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_6, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[18])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_90_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x3_sva_5, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[17])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_91_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_4, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[16])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_92_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_3, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[15])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_93_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_2, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[14])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_94_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_1, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[13])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_95_nl
      = MUX_s_1_2_2(rand_unit_random1_run_x2_12_0_sva_0, (~ (ac_math_atan_pi_2mi_return_2_69_28_sva[12])),
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_not_61_nl
      = ~ (fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_n000000
      = ~(MUX_v_12_2_2((ac_math_atan_pi_2mi_return_2_69_28_sva[11:0]), 12'b111111111111,
      (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_not_61_nl)));
  assign nl_acc_8_nl = conv_s2u_46_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_63_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_64_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_65_nl)
      , 1'b1}) + conv_s2u_45_47({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_if_or_1_cse
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_66_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_67_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_68_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_69_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_70_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_71_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_72_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_73_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_74_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_75_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_76_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_77_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_78_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_79_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_80_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_81_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_82_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_83_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_84_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_85_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_86_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_87_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_88_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_89_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_90_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_91_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_92_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_93_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_94_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_95_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_n000000)
      , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[46:0];
  assign z_out_8 = readslicef_47_46_1((acc_8_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_32_nl
      = MUX_v_3_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_44_42,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_33_nl
      = MUX_v_42_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_acc_a_lpi_1_dfm_1_41_0,
      fsm_output[13]);
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_34_nl
      = MUX_v_44_2_2(({lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21 ,
      lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_20_0 , 11'b00000000000}),
      ({2'b11 , (~ ac_math_atan_pi_2mi_return_69_28_sva)}), fsm_output[13]);
  assign nl_acc_9_nl = conv_s2u_46_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_32_nl)
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_33_nl)
      , 1'b1}) + conv_s2u_45_47({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_34_nl)
      , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[46:0];
  assign z_out_9 = readslicef_47_46_1((acc_9_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_nand_1_nl
      = ~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt
      & (~((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs)
      & (fsm_output[13]))));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_mux_29_nl
      = MUX_v_43_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_y_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_y_2mi_sva,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_9_rgt);
  assign nl_acc_10_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_35
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_32
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_18
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_15
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_x_lpi_1_dfm_1_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_nand_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_else_mux_29_nl)
      , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[43:0];
  assign z_out_10 = readslicef_44_43_1((acc_10_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_nand_1_nl
      = ~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt
      & (~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_slc_45_svs
      & (fsm_output[13]))));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_35_nl
      = MUX_v_43_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_x_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_x_2mi_sva,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_8_rgt);
  assign nl_acc_11_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_y_lpi_1_dfm_1_4_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_nand_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_for_if_mux_35_nl)
      , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[43:0];
  assign z_out_11 = readslicef_44_43_1((acc_11_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_1_nl
      = (~((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs)
      & (fsm_output[13]))) | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_29_nl
      = MUX_v_43_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_2mi_sva,
      (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_4_rgt);
  assign nl_acc_12_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_y_lpi_1_dfm_1_4_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_or_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_else_mux_29_nl)
      , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[43:0];
  assign z_out_12 = readslicef_44_43_1((acc_12_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_or_1_nl
      = (~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs
      & (fsm_output[13]))) | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_96_nl
      = MUX_v_43_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_y_2mi_sva,
      (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_y_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_7_cse);
  assign nl_acc_13_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_29
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_22
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_21
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_itm_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_x_lpi_1_dfm_1_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_or_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_if_mux_96_nl)
      , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[43:0];
  assign z_out_13 = readslicef_44_43_1((acc_13_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_nand_1_nl
      = ~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      & (~((~ ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_sel_lor_lpi_2_dfm_1)
      & (fsm_output[13]))));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_mux_29_nl
      = MUX_v_43_2_2((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_y_2mi_sva,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse);
  assign nl_acc_14_nl = ({ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_i_6_0_sva_1_3_0
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_2_itm_43_42
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_29
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_1_0
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_9
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_8
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_7
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_28
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_18_17
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_itm_15_14
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_22
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_20
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_16
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_x_lpi_1_dfm_1_5
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_x_d_acc_cse_7_0_sva_3_0
      , ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_mux_itm_12
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_nand_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_else_mux_29_nl)
      , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[43:0];
  assign z_out_14 = readslicef_44_43_1((acc_14_nl));
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_29_nl = MUX_v_4_2_2((signext_4_1(hit_in_crt_sva_171_0[140])),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_42_39,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_30_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_38,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_31_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_37,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_32_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_36,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_33_nl = MUX_v_2_2_2((signext_2_1(hit_in_crt_sva_171_0[140])),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_35_34,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_34_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_33,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_35_nl = MUX_v_2_2_2((signext_2_1(hit_in_crt_sva_171_0[140])),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_32_31,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_36_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_30,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_37_nl = MUX_v_3_2_2((signext_3_1(hit_in_crt_sva_171_0[140])),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_29_27,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_38_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_26,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_39_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[140]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_25,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_40_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[139]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_24,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_41_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[138]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_23,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_42_nl = MUX_v_3_2_2((hit_in_crt_sva_171_0[137:135]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_22_20,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_43_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[134]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_19,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_44_nl = MUX_v_2_2_2((hit_in_crt_sva_171_0[133:132]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_18_17,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_45_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[131]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_16,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_46_nl = MUX_v_2_2_2((hit_in_crt_sva_171_0[130:129]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_15_14,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_47_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[128]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_13,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_48_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[127]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_12,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_49_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[126]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_11,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_50_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[125]),
      ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_ac_math_ac_arccos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_acc_6_itm,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_51_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[124]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_9,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_52_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[123]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_8,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_53_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[122]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_7,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_54_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[121]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_6,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_55_nl = MUX_s_1_2_2((hit_in_crt_sva_171_0[120]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_mux_1_itm_5,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_56_nl = MUX_v_5_2_2((hit_in_crt_sva_171_0[119:115]),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_y_lpi_1_dfm_1_4_0,
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_or_16_rgt);
  assign lambertianScatter_add_run_or_30_nl = (~((fsm_output[14]) | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse))
      | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse;
  assign lambertianScatter_add_run_mux1h_44_nl = MUX1HOT_v_2_3_2((signext_2_1(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[25])),
      (~ reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd),
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd,
      {(fsm_output[14]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse});
  assign lambertianScatter_add_run_lambertianScatter_add_run_mux_57_nl = MUX_s_1_2_2((reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[25]),
      (~ (reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[25])),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse);
  assign lambertianScatter_add_run_mux1h_45_nl = MUX1HOT_v_25_3_2((signext_25_11(reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[25:15])),
      (~ (reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[24:0])),
      (reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[24:0]),
      {(fsm_output[14]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse});
  assign lambertianScatter_add_run_mux1h_46_nl = MUX1HOT_v_8_3_2((reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[14:7]),
      (~ reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2),
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_2,
      {(fsm_output[14]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse});
  assign lambertianScatter_add_run_mux1h_47_nl = MUX1HOT_v_7_3_2((reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_1[6:0]),
      (~ reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_3),
      reg_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_for_x_2mi_ftd_3,
      {(fsm_output[14]) , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_83_cse
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_and_82_cse});
  assign nl_acc_15_nl = ({(lambertianScatter_add_run_lambertianScatter_add_run_mux_29_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_30_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_31_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_32_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_33_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_34_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_35_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_36_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_37_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_38_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_39_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_40_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_41_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_42_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_43_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_44_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_45_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_46_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_47_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_48_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_49_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_50_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_51_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_52_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_53_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_54_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_55_nl)
      , (lambertianScatter_add_run_lambertianScatter_add_run_mux_56_nl) , (lambertianScatter_add_run_or_30_nl)})
      + ({(lambertianScatter_add_run_mux1h_44_nl) , (lambertianScatter_add_run_lambertianScatter_add_run_mux_57_nl)
      , (lambertianScatter_add_run_mux1h_45_nl) , (lambertianScatter_add_run_mux1h_46_nl)
      , (lambertianScatter_add_run_mux1h_47_nl) , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[43:0];
  assign z_out_15 = readslicef_44_43_1((acc_15_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_or_1_nl
      = (~((~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_slc_45_svs)
      & (fsm_output[13]))) | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_mux_29_nl
      = MUX_v_43_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_x_2mi_sva,
      (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_x_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_and_8_cse);
  assign nl_acc_16_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_37
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_35_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_32_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_24
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_18_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_15_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_9
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_8
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_7
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_mux_1_itm_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_y_lpi_1_dfm_1_4_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_or_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_2_for_else_mux_29_nl)
      , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[43:0];
  assign z_out_16 = readslicef_44_43_1((acc_16_nl));
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_or_1_nl
      = (~(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_slc_45_svs
      & (fsm_output[13]))) | ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_35_nl
      = MUX_v_43_2_2(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_sva,
      (~ ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_y_2mi_sva),
      ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_3_acc_a_and_3_rgt);
  assign nl_acc_17_nl = ({ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_42_39
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_38
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_37_36
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_35
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_34
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_33
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_32
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_31
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_30
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_29_27
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_26
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_25
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_24_23
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_22_20
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_19
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_18
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_17
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_16
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_15
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_14
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_13
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_12
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_11
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_10
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_9_6
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_5
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_4_1
      , ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_x_lpi_1_dfm_1_0
      , (ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_or_1_nl)})
      + ({(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_for_if_mux_35_nl)
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[43:0];
  assign z_out_17 = readslicef_44_43_1((acc_17_nl));
  assign lambertianScatter_add_run_mux_8_nl = MUX_v_26_2_2((lambertianScatter_run_aelse_1_slc_lambertianScatter_run_zz_33_6_itm_26_0[25:0]),
      color_out_g_sva_1_25_0, fsm_output[17]);
  assign nl_z_out_18 = conv_s2u_26_27(lambertianScatter_add_run_mux_8_nl) + conv_s2u_26_27(lambertianScatter_rand_unit_run_xs_mul_cmp_z_oreg[33:8]);
  assign z_out_18 = nl_z_out_18[26:0];
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_mux_1_nl
      = MUX_v_2_2_2(({rand_unit_random1_run_x3_sva_31 , rand_unit_random1_run_x3_sva_30}),
      (lambertianScatter_rand_unit_run_phi_32_0_lpi_1_dfm_32_21[11:10]), fsm_output[11]);
  assign nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl
      = conv_s2u_2_3(ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_mux_1_nl)
      + 3'b001;
  assign ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl
      = nl_ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl[2:0];
  assign z_out_21_2 = readslicef_3_1_2((ac_math_ac_sincos_cordic_36_4_AC_TRN_AC_WRAP_36_4_AC_TRN_AC_WRAP_1_else_if_acc_nl));

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [24:0] MUX1HOT_v_25_3_2;
    input [24:0] input_2;
    input [24:0] input_1;
    input [24:0] input_0;
    input [2:0] sel;
    reg [24:0] result;
  begin
    result = input_0 & {25{sel[0]}};
    result = result | ( input_1 & {25{sel[1]}});
    result = result | ( input_2 & {25{sel[2]}});
    MUX1HOT_v_25_3_2 = result;
  end
  endfunction


  function automatic [26:0] MUX1HOT_v_27_3_2;
    input [26:0] input_2;
    input [26:0] input_1;
    input [26:0] input_0;
    input [2:0] sel;
    reg [26:0] result;
  begin
    result = input_0 & {27{sel[0]}};
    result = result | ( input_1 & {27{sel[1]}});
    result = result | ( input_2 & {27{sel[2]}});
    MUX1HOT_v_27_3_2 = result;
  end
  endfunction


  function automatic [27:0] MUX1HOT_v_28_3_2;
    input [27:0] input_2;
    input [27:0] input_1;
    input [27:0] input_0;
    input [2:0] sel;
    reg [27:0] result;
  begin
    result = input_0 & {28{sel[0]}};
    result = result | ( input_1 & {28{sel[1]}});
    result = result | ( input_2 & {28{sel[2]}});
    MUX1HOT_v_28_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [32:0] MUX1HOT_v_33_3_2;
    input [32:0] input_2;
    input [32:0] input_1;
    input [32:0] input_0;
    input [2:0] sel;
    reg [32:0] result;
  begin
    result = input_0 & {33{sel[0]}};
    result = result | ( input_1 & {33{sel[1]}});
    result = result | ( input_2 & {33{sel[2]}});
    MUX1HOT_v_33_3_2 = result;
  end
  endfunction


  function automatic [35:0] MUX1HOT_v_36_4_2;
    input [35:0] input_3;
    input [35:0] input_2;
    input [35:0] input_1;
    input [35:0] input_0;
    input [3:0] sel;
    reg [35:0] result;
  begin
    result = input_0 & {36{sel[0]}};
    result = result | ( input_1 & {36{sel[1]}});
    result = result | ( input_2 & {36{sel[2]}});
    result = result | ( input_3 & {36{sel[3]}});
    MUX1HOT_v_36_4_2 = result;
  end
  endfunction


  function automatic [35:0] MUX1HOT_v_36_5_2;
    input [35:0] input_4;
    input [35:0] input_3;
    input [35:0] input_2;
    input [35:0] input_1;
    input [35:0] input_0;
    input [4:0] sel;
    reg [35:0] result;
  begin
    result = input_0 & {36{sel[0]}};
    result = result | ( input_1 & {36{sel[1]}});
    result = result | ( input_2 & {36{sel[2]}});
    result = result | ( input_3 & {36{sel[3]}});
    result = result | ( input_4 & {36{sel[4]}});
    MUX1HOT_v_36_5_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [65:0] MUX1HOT_v_66_3_2;
    input [65:0] input_2;
    input [65:0] input_1;
    input [65:0] input_0;
    input [2:0] sel;
    reg [65:0] result;
  begin
    result = input_0 & {66{sel[0]}};
    result = result | ( input_1 & {66{sel[1]}});
    result = result | ( input_2 & {66{sel[2]}});
    MUX1HOT_v_66_3_2 = result;
  end
  endfunction


  function automatic [68:0] MUX1HOT_v_69_3_2;
    input [68:0] input_2;
    input [68:0] input_1;
    input [68:0] input_0;
    input [2:0] sel;
    reg [68:0] result;
  begin
    result = input_0 & {69{sel[0]}};
    result = result | ( input_1 & {69{sel[1]}});
    result = result | ( input_2 & {69{sel[2]}});
    MUX1HOT_v_69_3_2 = result;
  end
  endfunction


  function automatic [68:0] MUX1HOT_v_69_4_2;
    input [68:0] input_3;
    input [68:0] input_2;
    input [68:0] input_1;
    input [68:0] input_0;
    input [3:0] sel;
    reg [68:0] result;
  begin
    result = input_0 & {69{sel[0]}};
    result = result | ( input_1 & {69{sel[1]}});
    result = result | ( input_2 & {69{sel[2]}});
    result = result | ( input_3 & {69{sel[3]}});
    MUX1HOT_v_69_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction


  function automatic [25:0] MUX_v_26_2_2;
    input [25:0] input_0;
    input [25:0] input_1;
    input [0:0] sel;
    reg [25:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_26_2_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_2_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input [0:0] sel;
    reg [26:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_27_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [33:0] MUX_v_34_2_2;
    input [33:0] input_0;
    input [33:0] input_1;
    input [0:0] sel;
    reg [33:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_34_2_2 = result;
  end
  endfunction


  function automatic [35:0] MUX_v_36_2_2;
    input [35:0] input_0;
    input [35:0] input_1;
    input [0:0] sel;
    reg [35:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_36_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [41:0] MUX_v_42_2_2;
    input [41:0] input_0;
    input [41:0] input_1;
    input [0:0] sel;
    reg [41:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_42_2_2 = result;
  end
  endfunction


  function automatic [41:0] MUX_v_42_37_2;
    input [41:0] input_0;
    input [41:0] input_1;
    input [41:0] input_2;
    input [41:0] input_3;
    input [41:0] input_4;
    input [41:0] input_5;
    input [41:0] input_6;
    input [41:0] input_7;
    input [41:0] input_8;
    input [41:0] input_9;
    input [41:0] input_10;
    input [41:0] input_11;
    input [41:0] input_12;
    input [41:0] input_13;
    input [41:0] input_14;
    input [41:0] input_15;
    input [41:0] input_16;
    input [41:0] input_17;
    input [41:0] input_18;
    input [41:0] input_19;
    input [41:0] input_20;
    input [41:0] input_21;
    input [41:0] input_22;
    input [41:0] input_23;
    input [41:0] input_24;
    input [41:0] input_25;
    input [41:0] input_26;
    input [41:0] input_27;
    input [41:0] input_28;
    input [41:0] input_29;
    input [41:0] input_30;
    input [41:0] input_31;
    input [41:0] input_32;
    input [41:0] input_33;
    input [41:0] input_34;
    input [41:0] input_35;
    input [41:0] input_36;
    input [5:0] sel;
    reg [41:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      default : begin
        result = input_36;
      end
    endcase
    MUX_v_42_37_2 = result;
  end
  endfunction


  function automatic [42:0] MUX_v_43_2_2;
    input [42:0] input_0;
    input [42:0] input_1;
    input [0:0] sel;
    reg [42:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_43_2_2 = result;
  end
  endfunction


  function automatic [43:0] MUX_v_44_2_2;
    input [43:0] input_0;
    input [43:0] input_1;
    input [0:0] sel;
    reg [43:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_44_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_66_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [63:0] input_2;
    input [63:0] input_3;
    input [63:0] input_4;
    input [63:0] input_5;
    input [63:0] input_6;
    input [63:0] input_7;
    input [63:0] input_8;
    input [63:0] input_9;
    input [63:0] input_10;
    input [63:0] input_11;
    input [63:0] input_12;
    input [63:0] input_13;
    input [63:0] input_14;
    input [63:0] input_15;
    input [63:0] input_16;
    input [63:0] input_17;
    input [63:0] input_18;
    input [63:0] input_19;
    input [63:0] input_20;
    input [63:0] input_21;
    input [63:0] input_22;
    input [63:0] input_23;
    input [63:0] input_24;
    input [63:0] input_25;
    input [63:0] input_26;
    input [63:0] input_27;
    input [63:0] input_28;
    input [63:0] input_29;
    input [63:0] input_30;
    input [63:0] input_31;
    input [63:0] input_32;
    input [63:0] input_33;
    input [63:0] input_34;
    input [63:0] input_35;
    input [63:0] input_36;
    input [63:0] input_37;
    input [63:0] input_38;
    input [63:0] input_39;
    input [63:0] input_40;
    input [63:0] input_41;
    input [63:0] input_42;
    input [63:0] input_43;
    input [63:0] input_44;
    input [63:0] input_45;
    input [63:0] input_46;
    input [63:0] input_47;
    input [63:0] input_48;
    input [63:0] input_49;
    input [63:0] input_50;
    input [63:0] input_51;
    input [63:0] input_52;
    input [63:0] input_53;
    input [63:0] input_54;
    input [63:0] input_55;
    input [63:0] input_56;
    input [63:0] input_57;
    input [63:0] input_58;
    input [63:0] input_59;
    input [63:0] input_60;
    input [63:0] input_61;
    input [63:0] input_62;
    input [63:0] input_63;
    input [63:0] input_64;
    input [63:0] input_65;
    input [6:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      default : begin
        result = input_65;
      end
    endcase
    MUX_v_64_66_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [65:0] MUX_v_66_2_2;
    input [65:0] input_0;
    input [65:0] input_1;
    input [0:0] sel;
    reg [65:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_66_2_2 = result;
  end
  endfunction


  function automatic [68:0] MUX_v_69_2_2;
    input [68:0] input_0;
    input [68:0] input_1;
    input [0:0] sel;
    reg [68:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_69_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [27:0] readslicef_34_28_6;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_34_28_6 = tmp[27:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [42:0] readslicef_44_43_1;
    input [43:0] vector;
    reg [43:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_44_43_1 = tmp[42:0];
  end
  endfunction


  function automatic [45:0] readslicef_47_46_1;
    input [46:0] vector;
    reg [46:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_47_46_1 = tmp[45:0];
  end
  endfunction


  function automatic [69:0] readslicef_71_70_1;
    input [70:0] vector;
    reg [70:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_71_70_1 = tmp[69:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [20:0] signext_21_1;
    input [0:0] vector;
  begin
    signext_21_1= {{20{vector[0]}}, vector};
  end
  endfunction


  function automatic [24:0] signext_25_11;
    input [10:0] vector;
  begin
    signext_25_11= {{14{vector[10]}}, vector};
  end
  endfunction


  function automatic [25:0] signext_26_1;
    input [0:0] vector;
  begin
    signext_26_1= {{25{vector[0]}}, vector};
  end
  endfunction


  function automatic [25:0] signext_26_25;
    input [24:0] vector;
  begin
    signext_26_25= {{1{vector[24]}}, vector};
  end
  endfunction


  function automatic [26:0] signext_27_1;
    input [0:0] vector;
  begin
    signext_27_1= {{26{vector[0]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [33:0] signext_34_1;
    input [0:0] vector;
  begin
    signext_34_1= {{33{vector[0]}}, vector};
  end
  endfunction


  function automatic [33:0] signext_34_26;
    input [25:0] vector;
  begin
    signext_34_26= {{8{vector[25]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function automatic [68:0] signext_69_43;
    input [42:0] vector;
  begin
    signext_69_43= {{26{vector[42]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_1;
    input [0:0] vector;
  begin
    signext_6_1= {{5{vector[0]}}, vector};
  end
  endfunction


  function automatic [65:0] conv_s2s_65_66 ;
    input [64:0]  vector ;
  begin
    conv_s2s_65_66 = {vector[64], vector};
  end
  endfunction


  function automatic [2:0] conv_s2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction


  function automatic [26:0] conv_s2u_26_27 ;
    input [25:0]  vector ;
  begin
    conv_s2u_26_27 = {vector[25], vector};
  end
  endfunction


  function automatic [33:0] conv_s2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_s2u_33_34 = {vector[32], vector};
  end
  endfunction


  function automatic [46:0] conv_s2u_45_47 ;
    input [44:0]  vector ;
  begin
    conv_s2u_45_47 = {{2{vector[44]}}, vector};
  end
  endfunction


  function automatic [46:0] conv_s2u_46_47 ;
    input [45:0]  vector ;
  begin
    conv_s2u_46_47 = {vector[45], vector};
  end
  endfunction


  function automatic [70:0] conv_s2u_70_71 ;
    input [69:0]  vector ;
  begin
    conv_s2u_70_71 = {vector[69], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [44:0] conv_u2s_42_45 ;
    input [41:0]  vector ;
  begin
    conv_u2s_42_45 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [65:0] conv_u2s_64_66 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_66 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_1_34 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_34 = {{33{1'b0}}, vector};
  end
  endfunction


  function automatic [28:0] conv_u2u_28_29 ;
    input [27:0]  vector ;
  begin
    conv_u2u_28_29 = {1'b0, vector};
  end
  endfunction


  function automatic [31:0] conv_u2u_31_32 ;
    input [30:0]  vector ;
  begin
    conv_u2u_31_32 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController_run
// ------------------------------------------------------------------


module ShaderFeedbackController_run (
  clk, arst_n, ray_chan_in_rsc_dat, ray_chan_in_rsc_vld, ray_chan_in_rsc_rdy, ray_scattered_chan_rsc_dat,
      ray_scattered_chan_rsc_vld, ray_scattered_chan_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, color_chan_in_rsc_dat, color_chan_in_rsc_vld,
      color_chan_in_rsc_rdy, atten_chan_in_rsc_dat, atten_chan_in_rsc_vld, atten_chan_in_rsc_rdy,
      ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, params_out_rsc_dat, params_out_rsc_vld,
      params_out_rsc_rdy, color_chan_out_rsc_dat, color_chan_out_rsc_vld, color_chan_out_rsc_rdy,
      atten_chan_out_rsc_dat, atten_chan_out_rsc_vld, atten_chan_out_rsc_rdy, output_pxl_serial_rsc_dat,
      output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_chan_in_rsc_dat;
  input ray_chan_in_rsc_vld;
  output ray_chan_in_rsc_rdy;
  input [165:0] ray_scattered_chan_rsc_dat;
  input ray_scattered_chan_rsc_vld;
  output ray_scattered_chan_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [80:0] color_chan_in_rsc_dat;
  input color_chan_in_rsc_vld;
  output color_chan_in_rsc_rdy;
  input [80:0] atten_chan_in_rsc_dat;
  input atten_chan_in_rsc_vld;
  output atten_chan_in_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;
  output [80:0] color_chan_out_rsc_dat;
  output color_chan_out_rsc_vld;
  input color_chan_out_rsc_rdy;
  output [80:0] atten_chan_out_rsc_dat;
  output atten_chan_out_rsc_vld;
  input atten_chan_out_rsc_rdy;
  output [80:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire ray_chan_in_rsci_wen_comp;
  wire [165:0] ray_chan_in_rsci_idat_mxwt;
  wire ray_scattered_chan_rsci_wen_comp;
  wire [165:0] ray_scattered_chan_rsci_idat_mxwt;
  wire params_in_rsci_wen_comp;
  wire [92:0] params_in_rsci_idat_mxwt;
  wire color_chan_in_rsci_wen_comp;
  wire [80:0] color_chan_in_rsci_idat_mxwt;
  wire atten_chan_in_rsci_wen_comp;
  wire [80:0] atten_chan_in_rsci_idat_mxwt;
  wire ray_out_rsci_wen_comp;
  wire params_out_rsci_wen_comp;
  reg [92:0] params_out_rsci_idat;
  wire color_chan_out_rsci_wen_comp;
  wire atten_chan_out_rsci_wen_comp;
  wire output_pxl_serial_rsci_wen_comp;
  reg [80:0] output_pxl_serial_rsci_idat;
  reg ray_out_rsci_idat_165;
  reg [33:0] ray_out_rsci_idat_164_131;
  reg [33:0] ray_out_rsci_idat_130_97;
  reg [33:0] ray_out_rsci_idat_96_63;
  reg [20:0] ray_out_rsci_idat_62_42;
  reg [20:0] ray_out_rsci_idat_41_21;
  reg [20:0] ray_out_rsci_idat_20_0;
  reg [26:0] color_chan_out_rsci_idat_80_54;
  reg [26:0] color_chan_out_rsci_idat_53_27;
  reg [26:0] color_chan_out_rsci_idat_26_0;
  reg [26:0] atten_chan_out_rsci_idat_80_54;
  reg [26:0] atten_chan_out_rsci_idat_53_27;
  reg [26:0] atten_chan_out_rsci_idat_26_0;
  wire [2:0] fsm_output;
  wire if_if_if_if_and_tmp;
  wire if_if_if_nand_tmp;
  wire or_tmp_1;
  wire atten_chan_out_and_cse;
  reg reg_output_pxl_serial_rsci_ivld_run_psct_cse;
  reg reg_atten_chan_out_rsci_ivld_run_psct_cse;
  reg reg_atten_chan_in_rsci_irdy_run_psct_cse;
  reg [1:0] iter_1_0_sva;
  reg [1:0] iter_3_2_sva;
  reg [32:0] sample_sva;
  wire [33:0] nl_sample_sva;
  wire [3:0] operator_4_false_acc_ncse_sva_1;
  wire [4:0] nl_operator_4_false_acc_ncse_sva_1;

  wire[0:0] oelse_not_7_nl;
  wire[0:0] oelse_not_4_nl;
  wire[0:0] oelse_not_6_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [165:0] nl_ShaderFeedbackController_run_ray_out_rsci_inst_ray_out_rsci_idat;
  assign nl_ShaderFeedbackController_run_ray_out_rsci_inst_ray_out_rsci_idat = {ray_out_rsci_idat_165
      , ray_out_rsci_idat_164_131 , ray_out_rsci_idat_130_97 , ray_out_rsci_idat_96_63
      , ray_out_rsci_idat_62_42 , ray_out_rsci_idat_41_21 , ray_out_rsci_idat_20_0};
  wire [80:0] nl_ShaderFeedbackController_run_color_chan_out_rsci_inst_color_chan_out_rsci_idat;
  assign nl_ShaderFeedbackController_run_color_chan_out_rsci_inst_color_chan_out_rsci_idat
      = {color_chan_out_rsci_idat_80_54 , color_chan_out_rsci_idat_53_27 , color_chan_out_rsci_idat_26_0};
  wire [80:0] nl_ShaderFeedbackController_run_atten_chan_out_rsci_inst_atten_chan_out_rsci_idat;
  assign nl_ShaderFeedbackController_run_atten_chan_out_rsci_inst_atten_chan_out_rsci_idat
      = {atten_chan_out_rsci_idat_80_54 , atten_chan_out_rsci_idat_53_27 , atten_chan_out_rsci_idat_26_0};
  ShaderFeedbackController_run_ray_chan_in_rsci ShaderFeedbackController_run_ray_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_chan_in_rsc_dat(ray_chan_in_rsc_dat),
      .ray_chan_in_rsc_vld(ray_chan_in_rsc_vld),
      .ray_chan_in_rsc_rdy(ray_chan_in_rsc_rdy),
      .run_wen(run_wen),
      .ray_chan_in_rsci_oswt(reg_atten_chan_in_rsci_irdy_run_psct_cse),
      .ray_chan_in_rsci_wen_comp(ray_chan_in_rsci_wen_comp),
      .ray_chan_in_rsci_idat_mxwt(ray_chan_in_rsci_idat_mxwt)
    );
  ShaderFeedbackController_run_ray_scattered_chan_rsci ShaderFeedbackController_run_ray_scattered_chan_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_scattered_chan_rsc_dat(ray_scattered_chan_rsc_dat),
      .ray_scattered_chan_rsc_vld(ray_scattered_chan_rsc_vld),
      .ray_scattered_chan_rsc_rdy(ray_scattered_chan_rsc_rdy),
      .run_wen(run_wen),
      .ray_scattered_chan_rsci_oswt(reg_atten_chan_in_rsci_irdy_run_psct_cse),
      .ray_scattered_chan_rsci_wen_comp(ray_scattered_chan_rsci_wen_comp),
      .ray_scattered_chan_rsci_idat_mxwt(ray_scattered_chan_rsci_idat_mxwt)
    );
  ShaderFeedbackController_run_params_in_rsci ShaderFeedbackController_run_params_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .run_wen(run_wen),
      .params_in_rsci_oswt(reg_atten_chan_in_rsci_irdy_run_psct_cse),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .params_in_rsci_idat_mxwt(params_in_rsci_idat_mxwt)
    );
  ShaderFeedbackController_run_color_chan_in_rsci ShaderFeedbackController_run_color_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .color_chan_in_rsc_dat(color_chan_in_rsc_dat),
      .color_chan_in_rsc_vld(color_chan_in_rsc_vld),
      .color_chan_in_rsc_rdy(color_chan_in_rsc_rdy),
      .run_wen(run_wen),
      .color_chan_in_rsci_oswt(reg_atten_chan_in_rsci_irdy_run_psct_cse),
      .color_chan_in_rsci_wen_comp(color_chan_in_rsci_wen_comp),
      .color_chan_in_rsci_idat_mxwt(color_chan_in_rsci_idat_mxwt)
    );
  ShaderFeedbackController_run_atten_chan_in_rsci ShaderFeedbackController_run_atten_chan_in_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .atten_chan_in_rsc_dat(atten_chan_in_rsc_dat),
      .atten_chan_in_rsc_vld(atten_chan_in_rsc_vld),
      .atten_chan_in_rsc_rdy(atten_chan_in_rsc_rdy),
      .run_wen(run_wen),
      .atten_chan_in_rsci_oswt(reg_atten_chan_in_rsci_irdy_run_psct_cse),
      .atten_chan_in_rsci_wen_comp(atten_chan_in_rsci_wen_comp),
      .atten_chan_in_rsci_idat_mxwt(atten_chan_in_rsci_idat_mxwt)
    );
  ShaderFeedbackController_run_ray_out_rsci ShaderFeedbackController_run_ray_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .run_wen(run_wen),
      .ray_out_rsci_oswt(reg_atten_chan_out_rsci_ivld_run_psct_cse),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .ray_out_rsci_idat(nl_ShaderFeedbackController_run_ray_out_rsci_inst_ray_out_rsci_idat[165:0])
    );
  ShaderFeedbackController_run_params_out_rsci ShaderFeedbackController_run_params_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .params_out_rsc_dat(params_out_rsc_dat),
      .params_out_rsc_vld(params_out_rsc_vld),
      .params_out_rsc_rdy(params_out_rsc_rdy),
      .run_wen(run_wen),
      .params_out_rsci_oswt(reg_atten_chan_out_rsci_ivld_run_psct_cse),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp),
      .params_out_rsci_idat(params_out_rsci_idat)
    );
  ShaderFeedbackController_run_color_chan_out_rsci ShaderFeedbackController_run_color_chan_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .color_chan_out_rsc_dat(color_chan_out_rsc_dat),
      .color_chan_out_rsc_vld(color_chan_out_rsc_vld),
      .color_chan_out_rsc_rdy(color_chan_out_rsc_rdy),
      .run_wen(run_wen),
      .color_chan_out_rsci_oswt(reg_atten_chan_out_rsci_ivld_run_psct_cse),
      .color_chan_out_rsci_wen_comp(color_chan_out_rsci_wen_comp),
      .color_chan_out_rsci_idat(nl_ShaderFeedbackController_run_color_chan_out_rsci_inst_color_chan_out_rsci_idat[80:0])
    );
  ShaderFeedbackController_run_atten_chan_out_rsci ShaderFeedbackController_run_atten_chan_out_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .atten_chan_out_rsc_dat(atten_chan_out_rsc_dat),
      .atten_chan_out_rsc_vld(atten_chan_out_rsc_vld),
      .atten_chan_out_rsc_rdy(atten_chan_out_rsc_rdy),
      .run_wen(run_wen),
      .atten_chan_out_rsci_oswt(reg_atten_chan_out_rsci_ivld_run_psct_cse),
      .atten_chan_out_rsci_wen_comp(atten_chan_out_rsci_wen_comp),
      .atten_chan_out_rsci_idat(nl_ShaderFeedbackController_run_atten_chan_out_rsci_inst_atten_chan_out_rsci_idat[80:0])
    );
  ShaderFeedbackController_run_output_pxl_serial_rsci ShaderFeedbackController_run_output_pxl_serial_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy),
      .run_wen(run_wen),
      .output_pxl_serial_rsci_oswt(reg_output_pxl_serial_rsci_ivld_run_psct_cse),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp),
      .output_pxl_serial_rsci_idat(output_pxl_serial_rsci_idat)
    );
  ShaderFeedbackController_run_staller ShaderFeedbackController_run_staller_inst
      (
      .run_wen(run_wen),
      .ray_chan_in_rsci_wen_comp(ray_chan_in_rsci_wen_comp),
      .ray_scattered_chan_rsci_wen_comp(ray_scattered_chan_rsci_wen_comp),
      .params_in_rsci_wen_comp(params_in_rsci_wen_comp),
      .color_chan_in_rsci_wen_comp(color_chan_in_rsci_wen_comp),
      .atten_chan_in_rsci_wen_comp(atten_chan_in_rsci_wen_comp),
      .ray_out_rsci_wen_comp(ray_out_rsci_wen_comp),
      .params_out_rsci_wen_comp(params_out_rsci_wen_comp),
      .color_chan_out_rsci_wen_comp(color_chan_out_rsci_wen_comp),
      .atten_chan_out_rsci_wen_comp(atten_chan_out_rsci_wen_comp),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp)
    );
  ShaderFeedbackController_run_run_fsm ShaderFeedbackController_run_run_fsm_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output)
    );
  assign atten_chan_out_and_cse = run_wen & (fsm_output[1]);
  assign if_if_if_nand_tmp = ~((~((iter_1_0_sva[0]) & (~((iter_3_2_sva!=2'b00) |
      (iter_1_0_sva[1]))))) & ((iter_3_2_sva!=2'b00) | (iter_1_0_sva!=2'b00)));
  assign nl_operator_4_false_acc_ncse_sva_1 = ({iter_3_2_sva , iter_1_0_sva}) + 4'b0001;
  assign operator_4_false_acc_ncse_sva_1 = nl_operator_4_false_acc_ncse_sva_1[3:0];
  assign if_if_if_if_and_tmp = (~((sample_sva[0]) & (~((sample_sva[32:4]!=29'b00000000000000000000000000000)))))
      & ((sample_sva[32]) | (sample_sva[31]) | (sample_sva[30]) | (sample_sva[29])
      | (sample_sva[28]) | (sample_sva[27]) | (sample_sva[26]) | (sample_sva[25])
      | (sample_sva[24]) | (sample_sva[23]) | (sample_sva[22]) | (sample_sva[21])
      | (sample_sva[20]) | (sample_sva[19]) | (sample_sva[18]) | (sample_sva[17])
      | (sample_sva[16]) | (sample_sva[15]) | (sample_sva[14]) | (sample_sva[13])
      | (sample_sva[12]) | (sample_sva[11]) | (sample_sva[10]) | (sample_sva[9])
      | (sample_sva[8]) | (sample_sva[7]) | (sample_sva[6]) | (sample_sva[5]) | (sample_sva[4])
      | (sample_sva[0]));
  assign or_tmp_1 = (~ if_if_if_nand_tmp) & (fsm_output[1]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      atten_chan_out_rsci_idat_26_0 <= 27'b000000000000000000000000000;
      atten_chan_out_rsci_idat_53_27 <= 27'b000000000000000000000000000;
      atten_chan_out_rsci_idat_80_54 <= 27'b000000000000000000000000000;
      color_chan_out_rsci_idat_26_0 <= 27'b000000000000000000000000000;
      color_chan_out_rsci_idat_53_27 <= 27'b000000000000000000000000000;
      color_chan_out_rsci_idat_80_54 <= 27'b000000000000000000000000000;
      ray_out_rsci_idat_20_0 <= 21'b000000000000000000000;
      ray_out_rsci_idat_41_21 <= 21'b000000000000000000000;
      ray_out_rsci_idat_62_42 <= 21'b000000000000000000000;
      ray_out_rsci_idat_96_63 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_130_97 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_164_131 <= 34'b0000000000000000000000000000000000;
      ray_out_rsci_idat_165 <= 1'b0;
      params_out_rsci_idat <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      sample_sva <= 33'b000000000000000000000000000000000;
      iter_1_0_sva <= 2'b00;
      iter_3_2_sva <= 2'b00;
    end
    else if ( atten_chan_out_and_cse ) begin
      atten_chan_out_rsci_idat_26_0 <= MUX_v_27_2_2(27'b000010000000000000000000000,
          (atten_chan_in_rsci_idat_mxwt[26:0]), or_tmp_1);
      atten_chan_out_rsci_idat_53_27 <= MUX_v_27_2_2(27'b000010000000000000000000000,
          (atten_chan_in_rsci_idat_mxwt[53:27]), or_tmp_1);
      atten_chan_out_rsci_idat_80_54 <= MUX_v_27_2_2(27'b000010000000000000000000000,
          (atten_chan_in_rsci_idat_mxwt[80:54]), or_tmp_1);
      color_chan_out_rsci_idat_26_0 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (color_chan_in_rsci_idat_mxwt[26:0]), (oelse_not_7_nl));
      color_chan_out_rsci_idat_53_27 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (color_chan_in_rsci_idat_mxwt[53:27]), (oelse_not_4_nl));
      color_chan_out_rsci_idat_80_54 <= MUX_v_27_2_2(27'b000000000000000000000000000,
          (color_chan_in_rsci_idat_mxwt[80:54]), (oelse_not_6_nl));
      ray_out_rsci_idat_20_0 <= MUX_v_21_2_2((ray_chan_in_rsci_idat_mxwt[20:0]),
          (ray_scattered_chan_rsci_idat_mxwt[20:0]), or_tmp_1);
      ray_out_rsci_idat_41_21 <= MUX_v_21_2_2((ray_chan_in_rsci_idat_mxwt[41:21]),
          (ray_scattered_chan_rsci_idat_mxwt[41:21]), or_tmp_1);
      ray_out_rsci_idat_62_42 <= MUX_v_21_2_2((ray_chan_in_rsci_idat_mxwt[62:42]),
          (ray_scattered_chan_rsci_idat_mxwt[62:42]), or_tmp_1);
      ray_out_rsci_idat_96_63 <= MUX_v_34_2_2((ray_chan_in_rsci_idat_mxwt[96:63]),
          (ray_scattered_chan_rsci_idat_mxwt[96:63]), or_tmp_1);
      ray_out_rsci_idat_130_97 <= MUX_v_34_2_2((ray_chan_in_rsci_idat_mxwt[130:97]),
          (ray_scattered_chan_rsci_idat_mxwt[130:97]), or_tmp_1);
      ray_out_rsci_idat_164_131 <= MUX_v_34_2_2((ray_chan_in_rsci_idat_mxwt[164:131]),
          (ray_scattered_chan_rsci_idat_mxwt[164:131]), or_tmp_1);
      ray_out_rsci_idat_165 <= MUX_s_1_2_2((ray_chan_in_rsci_idat_mxwt[165]), (ray_scattered_chan_rsci_idat_mxwt[165]),
          or_tmp_1);
      params_out_rsci_idat <= params_in_rsci_idat_mxwt;
      sample_sva <= nl_sample_sva[32:0];
      iter_1_0_sva <= operator_4_false_acc_ncse_sva_1[1:0];
      iter_3_2_sva <= operator_4_false_acc_ncse_sva_1[3:2];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_pxl_serial_rsci_idat <= 81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( run_wen & if_if_if_nand_tmp & if_if_if_if_and_tmp & (fsm_output[1])
        ) begin
      output_pxl_serial_rsci_idat <= color_chan_in_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_output_pxl_serial_rsci_ivld_run_psct_cse <= 1'b0;
      reg_atten_chan_out_rsci_ivld_run_psct_cse <= 1'b0;
      reg_atten_chan_in_rsci_irdy_run_psct_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_output_pxl_serial_rsci_ivld_run_psct_cse <= if_if_if_nand_tmp & if_if_if_if_and_tmp
          & (fsm_output[1]);
      reg_atten_chan_out_rsci_ivld_run_psct_cse <= fsm_output[1];
      reg_atten_chan_in_rsci_irdy_run_psct_cse <= ~ (fsm_output[1]);
    end
  end
  assign oelse_not_7_nl = ~ if_if_if_nand_tmp;
  assign oelse_not_4_nl = ~ if_if_if_nand_tmp;
  assign oelse_not_6_nl = ~ if_if_if_nand_tmp;
  assign nl_sample_sva  = sample_sva + 33'b000000000000000000000000000000001;

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction


  function automatic [26:0] MUX_v_27_2_2;
    input [26:0] input_0;
    input [26:0] input_1;
    input [0:0] sel;
    reg [26:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_27_2_2 = result;
  end
  endfunction


  function automatic [33:0] MUX_v_34_2_2;
    input [33:0] input_0;
    input [33:0] input_1;
    input [0:0] sel;
    reg [33:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_34_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector_run
// ------------------------------------------------------------------


module RayCollector_run (
  clk, arst_n, rayIn_rsc_dat, rayIn_rsc_vld, rayIn_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy,
      rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] rayIn_rsc_dat;
  input rayIn_rsc_vld;
  output rayIn_rsc_rdy;
  input [92:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire rayIn_rsci_wen_comp;
  wire [165:0] rayIn_rsci_idat_mxwt;
  wire paramsIn_rsci_wen_comp;
  wire [92:0] paramsIn_rsci_idat_mxwt;
  wire paramsOut_rsci_wen_comp;
  reg [92:0] paramsOut_rsci_idat;
  wire rayOut_rsci_wen_comp;
  reg [165:0] rayOut_rsci_idat;
  wire [5:0] fsm_output;
  wire and_21_cse;
  reg for_slc_for_acc_4_itm;
  reg [92:0] paramsIn_crt_1_sva;
  reg for_if_for_if_or_itm;
  reg [3:0] for_i_3_0_sva;
  reg reg_rayOut_rsci_ivld_run_psct_cse;
  wire rayOut_and_cse;
  reg reg_paramsIn_rsci_irdy_run_psct_cse;
  wire for_if_for_if_or_cse;
  wire rayOut_or_itm;
  reg [92:0] paramsIn_crt_sva;
  reg [165:0] rayIn_crt_sva;
  reg [165:0] rayIn_crt_1_sva;
  wire [3:0] for_i_3_0_sva_1_mx0w1;
  wire [4:0] nl_for_i_3_0_sva_1_mx0w1;
  wire and_cse;
  wire and_55_cse;

  wire[0:0] nor_2_nl;
  wire[4:0] for_acc_nl;
  wire[5:0] nl_for_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_RayCollector_run_run_fsm_inst_for_C_2_tr0;
  assign nl_RayCollector_run_run_fsm_inst_for_C_2_tr0 = ~ for_slc_for_acc_4_itm;
  RayCollector_run_rayIn_rsci RayCollector_run_rayIn_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rayIn_rsc_dat(rayIn_rsc_dat),
      .rayIn_rsc_vld(rayIn_rsc_vld),
      .rayIn_rsc_rdy(rayIn_rsc_rdy),
      .run_wen(run_wen),
      .rayIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .rayIn_rsci_wen_comp(rayIn_rsci_wen_comp),
      .rayIn_rsci_idat_mxwt(rayIn_rsci_idat_mxwt)
    );
  RayCollector_run_paramsIn_rsci RayCollector_run_paramsIn_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .run_wen(run_wen),
      .paramsIn_rsci_oswt(reg_paramsIn_rsci_irdy_run_psct_cse),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsIn_rsci_idat_mxwt(paramsIn_rsci_idat_mxwt)
    );
  RayCollector_run_paramsOut_rsci RayCollector_run_paramsOut_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .run_wen(run_wen),
      .paramsOut_rsci_oswt(reg_rayOut_rsci_ivld_run_psct_cse),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .paramsOut_rsci_idat(paramsOut_rsci_idat)
    );
  RayCollector_run_rayOut_rsci RayCollector_run_rayOut_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rayOut_rsc_dat(rayOut_rsc_dat),
      .rayOut_rsc_vld(rayOut_rsc_vld),
      .rayOut_rsc_rdy(rayOut_rsc_rdy),
      .run_wen(run_wen),
      .rayOut_rsci_oswt(reg_rayOut_rsci_ivld_run_psct_cse),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp),
      .rayOut_rsci_idat(rayOut_rsci_idat)
    );
  RayCollector_run_staller RayCollector_run_staller_inst (
      .run_wen(run_wen),
      .rayIn_rsci_wen_comp(rayIn_rsci_wen_comp),
      .paramsIn_rsci_wen_comp(paramsIn_rsci_wen_comp),
      .paramsOut_rsci_wen_comp(paramsOut_rsci_wen_comp),
      .rayOut_rsci_wen_comp(rayOut_rsci_wen_comp)
    );
  RayCollector_run_run_fsm RayCollector_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_C_2_tr0(nl_RayCollector_run_run_fsm_inst_for_C_2_tr0[0:0])
    );
  assign rayOut_or_itm = (for_if_for_if_or_cse & (fsm_output[3])) | and_21_cse;
  assign rayOut_and_cse = run_wen & rayOut_or_itm;
  assign and_cse = run_wen & ((fsm_output[1:0]!=2'b00));
  assign and_55_cse = run_wen & (fsm_output[5:3]==3'b000);
  assign for_if_for_if_or_cse = (paramsIn_crt_1_sva[92]) | (~ (for_i_3_0_sva[3]));
  assign nl_for_i_3_0_sva_1_mx0w1 = for_i_3_0_sva + 4'b0001;
  assign for_i_3_0_sva_1_mx0w1 = nl_for_i_3_0_sva_1_mx0w1[3:0];
  assign and_21_cse = for_if_for_if_or_itm & (fsm_output[4]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayOut_rsci_idat <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      paramsOut_rsci_idat <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( rayOut_and_cse ) begin
      rayOut_rsci_idat <= MUX_v_166_2_2(rayIn_crt_sva, rayIn_crt_1_sva, and_21_cse);
      paramsOut_rsci_idat <= MUX_v_93_2_2(paramsIn_crt_sva, paramsIn_crt_1_sva, and_21_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_rayOut_rsci_ivld_run_psct_cse <= 1'b0;
      reg_paramsIn_rsci_irdy_run_psct_cse <= 1'b0;
      for_if_for_if_or_itm <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_rayOut_rsci_ivld_run_psct_cse <= rayOut_or_itm;
      reg_paramsIn_rsci_irdy_run_psct_cse <= ~((fsm_output[4:2]!=3'b000) | (for_slc_for_acc_4_itm
          & (fsm_output[5])));
      for_if_for_if_or_itm <= for_if_for_if_or_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayIn_crt_sva <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      paramsIn_crt_sva <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_cse ) begin
      rayIn_crt_sva <= rayIn_rsci_idat_mxwt;
      paramsIn_crt_sva <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      rayIn_crt_1_sva <= 166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      paramsIn_crt_1_sva <= 93'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_55_cse ) begin
      rayIn_crt_1_sva <= rayIn_rsci_idat_mxwt;
      paramsIn_crt_1_sva <= paramsIn_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_i_3_0_sva <= 4'b0000;
    end
    else if ( (fsm_output[5:4]==2'b00) & run_wen ) begin
      for_i_3_0_sva <= MUX_v_4_2_2(4'b0000, for_i_3_0_sva_1_mx0w1, (nor_2_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_slc_for_acc_4_itm <= 1'b0;
    end
    else if ( run_wen & (fsm_output[3]) ) begin
      for_slc_for_acc_4_itm <= readslicef_5_1_4((for_acc_nl));
    end
  end
  assign nor_2_nl = ~((fsm_output[2:0]!=3'b000));
  assign nl_for_acc_nl = conv_u2s_4_5(for_i_3_0_sva_1_mx0w1) + 5'b10111;
  assign for_acc_nl = nl_for_acc_nl[4:0];

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [92:0] MUX_v_93_2_2;
    input [92:0] input_0;
    input [92:0] input_1;
    input [0:0] sel;
    reg [92:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_93_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator_run
// ------------------------------------------------------------------


module PixelAccumulator_run (
  clk, arst_n, accumulator_parms_rsc_dat, accumulator_parms_rsc_vld, accumulator_parms_rsc_rdy,
      pxl_sample_rsc_dat, pxl_sample_rsc_vld, pxl_sample_rsc_rdy, output_pxl_serial_rsc_dat,
      output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [419:0] accumulator_parms_rsc_dat;
  input accumulator_parms_rsc_vld;
  output accumulator_parms_rsc_rdy;
  input [80:0] pxl_sample_rsc_dat;
  input pxl_sample_rsc_vld;
  output pxl_sample_rsc_rdy;
  output [23:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire accumulator_parms_rsci_wen_comp;
  wire [34:0] accumulator_parms_rsci_idat_mxwt;
  wire pxl_sample_rsci_wen_comp;
  wire [80:0] pxl_sample_rsci_idat_mxwt;
  wire output_pxl_serial_rsci_wen_comp;
  reg output_pxl_serial_rsci_idat_23;
  reg output_pxl_serial_rsci_idat_22;
  reg output_pxl_serial_rsci_idat_21;
  reg output_pxl_serial_rsci_idat_20;
  reg output_pxl_serial_rsci_idat_19;
  reg output_pxl_serial_rsci_idat_18;
  reg output_pxl_serial_rsci_idat_17;
  reg output_pxl_serial_rsci_idat_16;
  reg output_pxl_serial_rsci_idat_15;
  reg output_pxl_serial_rsci_idat_14;
  reg output_pxl_serial_rsci_idat_13;
  reg output_pxl_serial_rsci_idat_12;
  reg output_pxl_serial_rsci_idat_11;
  reg output_pxl_serial_rsci_idat_10;
  reg output_pxl_serial_rsci_idat_9;
  reg output_pxl_serial_rsci_idat_8;
  reg output_pxl_serial_rsci_idat_7;
  reg output_pxl_serial_rsci_idat_6;
  reg output_pxl_serial_rsci_idat_5;
  reg output_pxl_serial_rsci_idat_4;
  reg output_pxl_serial_rsci_idat_3;
  reg output_pxl_serial_rsci_idat_2;
  reg output_pxl_serial_rsci_idat_1;
  reg output_pxl_serial_rsci_idat_0;
  wire [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_239_tmp;
  wire [11:0] for_acc_2_tmp;
  wire [12:0] nl_for_acc_2_tmp;
  wire operator_11_false_1_equal_1_tmp;
  wire [11:0] for_for_acc_1_tmp;
  wire [12:0] nl_for_for_acc_1_tmp;
  wire operator_11_false_equal_tmp;
  wire [4:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp;
  wire [5:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp;
  wire [4:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp;
  wire [5:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp;
  wire [4:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp;
  wire [5:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp;
  wire [1:0] for_mux_tmp;
  wire [16:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp;
  wire [18:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp;
  wire [16:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp;
  wire [18:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp;
  wire [16:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp;
  wire [18:0] nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp;
  wire or_tmp_7;
  wire or_dcpl_2;
  wire or_dcpl_4;
  wire and_dcpl_7;
  wire lfst_exit_for_for_lpi_1_dfm_mx0;
  wire exitL_exit_for_sva_mx0;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1;
  wire exit_for_for_for_lpi_1_dfm_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  wire exit_for_for_lpi_1_dfm_3;
  reg [1:0] lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_37_cse_1;
  reg [9:0] for_for_for_samps_10_0_lpi_1_dfm_1_9_0;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_23_cse_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_36_cse_1;
  wire for_for_else_3_unequal_tmp_1;
  wire for_for_for_unequal_tmp_1;
  wire for_for_blue_of_lpi_1_dfm_7_mx0;
  reg for_for_blue_of_lpi_1_dfm_1;
  wire for_for_green_of_lpi_1_dfm_7_mx0;
  reg for_for_green_of_lpi_1_dfm_1;
  wire for_for_red_of_lpi_1_dfm_7_mx0;
  reg for_for_red_of_lpi_1_dfm_1;
  wire for_for_for_and_2_tmp_1;
  wire for_for_for_and_1_tmp_1;
  wire for_for_for_and_tmp_1;
  reg exitL_exit_for_sva;
  reg main_stage_0_2;
  wire exit_for_lpi_1_dfm_3_mx0w0;
  reg exit_for_sva_2;
  wire [10:0] for_for_for_samps_10_0_sva_2;
  wire [11:0] nl_for_for_for_samps_10_0_sva_2;
  wire exit_for_for_for_sva_1;
  wire [6:0] operator_11_false_1_acc_sdt_sva_1;
  wire [7:0] nl_operator_11_false_1_acc_sdt_sva_1;
  wire [32:0] for_for_for_ac_fixed_cctor_2_sva_1;
  wire [33:0] nl_for_for_for_ac_fixed_cctor_2_sva_1;
  wire [32:0] for_for_for_ac_fixed_cctor_1_sva_1;
  wire [33:0] nl_for_for_for_ac_fixed_cctor_1_sva_1;
  wire [32:0] for_for_for_ac_fixed_cctor_sva_1;
  wire [33:0] nl_for_for_for_ac_fixed_cctor_sva_1;
  wire accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_94_cse_1;
  wire [1:0] lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_3;
  wire accumulator_parms_crt_lpi_1_dfm_12_11_mx2_1;
  wire [1:0] lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_4;
  reg reg_accumulator_parms_rsci_oswt_cse;
  reg reg_output_pxl_serial_rsci_oswt_cse;
  wire output_pxl_serial_and_cse;
  reg reg_pxl_sample_rsci_oswt_cse;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_and_cse;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_and_2_cse;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_and_cse;
  wire or_20_cse;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_9_8_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_7_6_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_11_10_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_5_4_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_13_12_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_3_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_14_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_1_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_9_8_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_7_6_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_11_10_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_5_4_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_13_12_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_3_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_14_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_1_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_9_8_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_7_6_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_11_10_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_5_4_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_13_12_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_3_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_14_lpi_1;
  reg [1:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_1_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_0_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_14_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
  reg ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1;
  reg [10:0] operator_12_true_return_10_0_lpi_1_dfm;
  reg [10:0] operator_11_false_return_10_0_lpi_1_dfm;
  reg mgc_qr_10_lpi_1_dfm_1;
  reg mgc_qr_8_lpi_1_dfm_1;
  reg mgc_qr_6_lpi_1_dfm_1;
  reg operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm;
  reg exit_for_for_for_sva;
  reg [32:0] for_for_accumulation_reg_x_lpi_1_dfm_1;
  reg [32:0] for_for_accumulation_reg_y_lpi_1_dfm_1;
  reg [32:0] for_for_accumulation_reg_z_lpi_1_dfm_1;
  reg [3:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_i_4_0_lpi_1_3_0;
  reg [3:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_i_4_0_lpi_1_3_0;
  reg [3:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_4_0_lpi_1_3_0;
  reg [1:0] accumulator_parms_crt_lpi_1_dfm_12_11;
  reg [10:0] for_fy_11_0_lpi_1_dfm_1_10_0;
  reg [10:0] for_for_fx_11_0_lpi_1_dfm_1_10_0;
  wire operator_2_false_2_operator_2_false_2_and_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_and_mdf_sva_1;
  wire operator_2_false_operator_2_false_nor_mdf_sva_1;
  wire mgc_qr_10_lpi_1_dfm_1_mx0;
  wire mgc_qr_8_lpi_1_dfm_1_mx0;
  wire mgc_qr_6_lpi_1_dfm_1_mx0;
  wire operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm_mx0;
  wire [10:0] operator_12_true_return_10_0_lpi_1_dfm_mx0;
  wire [10:0] operator_11_false_return_10_0_lpi_1_dfm_mx0;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_12_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_11_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_10_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_9_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_8_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_7_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_6_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_5_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_4_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_3_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_2_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_1_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_0_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_12_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_11_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_10_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_9_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_8_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_7_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_6_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_5_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_4_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_3_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_2_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_1_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_0_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_12_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_11_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_10_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_9_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_8_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_7_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_6_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_5_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_4_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_3_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_2_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_1_sva_1;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_0_sva_1;
  wire [14:0] for_for_rounded_accuracy_col_z_lpi_1_dfm_3;
  wire [14:0] for_for_rounded_accuracy_col_y_lpi_1_dfm_3;
  wire [14:0] for_for_rounded_accuracy_col_x_lpi_1_dfm_3;
  wire [19:0] for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1;
  wire [19:0] for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1;
  wire [19:0] for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1;
  wire for_for_asn_17;
  wire for_for_asn_19;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490;
  wire ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492;
  wire operator_33_true_equal_tmp;
  wire nand_3_cse;
  wire nor_8_cse;
  wire nor_23_cse;
  wire and_69_cse;
  wire and_81_cse;
  wire and_27_cse;

  wire[0:0] nor_nl;
  wire[9:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_96_nl;
  wire[0:0] mux_nl;
  wire[0:0] nand_14_nl;
  wire[0:0] and_89_nl;
  wire[0:0] for_not_20_nl;
  wire[10:0] for_for_for_for_for_for_mux_nl;
  wire[0:0] for_for_and_9_nl;
  wire[0:0] for_for_for_for_not_nl;
  wire[0:0] for_for_for_for_for_for_and_77_nl;
  wire[0:0] for_for_for_for_for_for_and_76_nl;
  wire[0:0] for_for_for_for_for_for_and_24_nl;
  wire[0:0] for_for_for_for_for_for_and_16_nl;
  wire[0:0] for_for_for_for_for_for_and_78_nl;
  wire[0:0] for_for_for_for_for_for_and_23_nl;
  wire[0:0] for_for_for_for_for_for_and_79_nl;
  wire[0:0] for_for_for_for_for_for_and_22_nl;
  wire[0:0] for_for_for_for_for_for_and_80_nl;
  wire[0:0] for_for_for_for_for_for_and_21_nl;
  wire[0:0] for_for_for_for_for_for_and_81_nl;
  wire[0:0] for_for_for_for_for_for_and_20_nl;
  wire[0:0] for_for_for_for_for_for_and_82_nl;
  wire[0:0] for_for_for_for_for_for_and_19_nl;
  wire[0:0] for_for_for_for_for_for_and_83_nl;
  wire[0:0] for_for_for_for_for_for_and_18_nl;
  wire[0:0] for_for_for_for_for_for_and_84_nl;
  wire[0:0] for_for_for_for_for_for_and_17_nl;
  wire[0:0] for_for_for_for_for_for_and_47_nl;
  wire[0:0] for_for_for_for_for_for_and_46_nl;
  wire[0:0] for_for_for_for_for_for_and_54_nl;
  wire[0:0] for_for_for_for_for_for_and_48_nl;
  wire[0:0] for_for_for_for_for_for_and_53_nl;
  wire[0:0] for_for_for_for_for_for_and_49_nl;
  wire[0:0] for_for_for_for_for_for_and_52_nl;
  wire[0:0] for_for_for_for_for_for_and_50_nl;
  wire[0:0] for_for_for_for_for_for_and_51_nl;
  wire[0:0] for_for_for_for_for_for_and_85_nl;
  wire[0:0] for_for_for_for_for_for_and_55_nl;
  wire[0:0] for_for_for_for_for_for_and_25_nl;
  wire[0:0] for_for_for_for_for_for_and_86_nl;
  wire[0:0] for_for_for_for_for_for_and_56_nl;
  wire[0:0] for_for_for_for_for_for_and_26_nl;
  wire[0:0] for_for_for_for_for_for_and_87_nl;
  wire[0:0] for_for_for_for_for_for_and_57_nl;
  wire[0:0] for_for_for_for_for_for_and_27_nl;
  wire[0:0] for_for_for_for_for_for_and_88_nl;
  wire[0:0] for_for_for_for_for_for_and_58_nl;
  wire[0:0] for_for_for_for_for_for_and_28_nl;
  wire[0:0] for_for_for_for_for_for_and_89_nl;
  wire[0:0] for_for_for_for_for_for_and_59_nl;
  wire[0:0] for_for_for_for_for_for_and_29_nl;
  wire[0:0] for_for_for_for_for_for_and_106_nl;
  wire[0:0] for_for_for_for_for_for_and_61_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_14_nl;
  wire[0:0] for_for_for_for_for_for_and_107_nl;
  wire[0:0] for_for_for_for_for_for_and_62_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_12_nl;
  wire[0:0] for_for_for_for_for_for_and_60_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_65_nl;
  wire[0:0] for_for_for_for_for_for_and_113_nl;
  wire[0:0] for_for_for_for_for_for_and_75_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_2_nl;
  wire[0:0] for_for_for_for_for_for_and_74_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_3_nl;
  wire[0:0] for_for_for_for_for_for_and_63_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_10_nl;
  wire[0:0] for_for_for_for_for_for_and_112_nl;
  wire[0:0] for_for_for_for_for_for_and_73_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_9_nl;
  wire[0:0] for_for_for_for_for_for_and_108_nl;
  wire[0:0] for_for_for_for_for_for_and_64_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_8_nl;
  wire[0:0] for_for_for_for_for_for_and_72_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_7_nl;
  wire[0:0] for_for_for_for_for_for_and_65_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_6_nl;
  wire[0:0] for_for_for_for_for_for_and_111_nl;
  wire[0:0] for_for_for_for_for_for_and_71_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_5_nl;
  wire[0:0] for_for_for_for_for_for_and_109_nl;
  wire[0:0] for_for_for_for_for_for_and_66_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_4_nl;
  wire[0:0] for_for_for_for_for_for_and_70_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_3_nl;
  wire[0:0] for_for_for_for_for_for_and_67_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_2_nl;
  wire[0:0] for_for_for_for_for_for_and_110_nl;
  wire[0:0] for_for_for_for_for_for_and_69_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_1_nl;
  wire[0:0] for_for_for_for_for_for_and_68_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_nl;
  wire[0:0] for_for_for_for_for_for_and_98_nl;
  wire[0:0] for_for_for_for_for_for_and_31_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_14_nl;
  wire[0:0] for_for_for_for_for_for_and_99_nl;
  wire[0:0] for_for_for_for_for_for_and_32_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_12_nl;
  wire[0:0] for_for_for_for_for_for_and_30_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_64_nl;
  wire[0:0] for_for_for_for_for_for_and_105_nl;
  wire[0:0] for_for_for_for_for_for_and_45_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_2_nl;
  wire[0:0] for_for_for_for_for_for_and_44_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_3_nl;
  wire[0:0] for_for_for_for_for_for_and_33_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_10_nl;
  wire[0:0] for_for_for_for_for_for_and_104_nl;
  wire[0:0] for_for_for_for_for_for_and_43_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_9_nl;
  wire[0:0] for_for_for_for_for_for_and_100_nl;
  wire[0:0] for_for_for_for_for_for_and_34_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_8_nl;
  wire[0:0] for_for_for_for_for_for_and_42_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_7_nl;
  wire[0:0] for_for_for_for_for_for_and_35_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_6_nl;
  wire[0:0] for_for_for_for_for_for_and_103_nl;
  wire[0:0] for_for_for_for_for_for_and_41_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_5_nl;
  wire[0:0] for_for_for_for_for_for_and_101_nl;
  wire[0:0] for_for_for_for_for_for_and_36_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_4_nl;
  wire[0:0] for_for_for_for_for_for_and_40_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_3_nl;
  wire[0:0] for_for_for_for_for_for_and_37_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_2_nl;
  wire[0:0] for_for_for_for_for_for_and_102_nl;
  wire[0:0] for_for_for_for_for_for_and_39_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_1_nl;
  wire[0:0] for_for_for_for_for_for_and_38_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_nl;
  wire[0:0] for_for_for_for_for_for_and_90_nl;
  wire[0:0] for_for_for_for_for_for_and_1_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_14_nl;
  wire[0:0] for_for_for_for_for_for_and_91_nl;
  wire[0:0] for_for_for_for_for_for_and_2_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_12_nl;
  wire[0:0] for_for_for_for_for_for_and_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_63_nl;
  wire[0:0] for_for_for_for_for_for_and_97_nl;
  wire[0:0] for_for_for_for_for_for_and_15_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_2_nl;
  wire[0:0] for_for_for_for_for_for_and_14_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_3_nl;
  wire[0:0] for_for_for_for_for_for_and_3_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_10_nl;
  wire[0:0] for_for_for_for_for_for_and_96_nl;
  wire[0:0] for_for_for_for_for_for_and_13_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_9_nl;
  wire[0:0] for_for_for_for_for_for_and_92_nl;
  wire[0:0] for_for_for_for_for_for_and_4_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_8_nl;
  wire[0:0] for_for_for_for_for_for_and_12_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_7_nl;
  wire[0:0] for_for_for_for_for_for_and_5_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_6_nl;
  wire[0:0] for_for_for_for_for_for_and_95_nl;
  wire[0:0] for_for_for_for_for_for_and_11_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_5_nl;
  wire[0:0] for_for_for_for_for_for_and_93_nl;
  wire[0:0] for_for_for_for_for_for_and_6_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_4_nl;
  wire[0:0] for_for_for_for_for_for_and_10_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_3_nl;
  wire[0:0] for_for_for_for_for_for_and_7_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_2_nl;
  wire[0:0] for_for_for_for_for_for_and_94_nl;
  wire[0:0] for_for_for_for_for_for_and_9_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_1_nl;
  wire[0:0] for_for_for_for_for_for_and_8_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_5_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_10_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_4_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_9_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_3_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_8_nl;
  wire[32:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_2_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_172_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_173_nl;
  wire[32:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_1_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_170_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_171_nl;
  wire[32:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_168_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_169_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] nor_12_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_174_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_175_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_37_nl;
  wire[0:0] for_mux_6_nl;
  wire[0:0] nor_1_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_nl;
  wire[10:0] operator_12_true_acc_nl;
  wire[11:0] nl_operator_12_true_acc_nl;
  wire[10:0] operator_11_false_acc_nl;
  wire[11:0] nl_operator_11_false_acc_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_14_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_12_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_14_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_12_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_14_nl;
  wire[0:0] ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_12_nl;
  wire[0:0] for_for_for_else_mux_3_nl;
  wire[0:0] for_for_for_else_if_for_for_for_else_if_or_2_nl;
  wire[0:0] for_for_for_else_else_mux_2_nl;
  wire[0:0] for_for_for_else_else_else_for_for_for_else_else_else_or_2_nl;
  wire[0:0] for_for_for_else_else_if_for_for_for_else_else_if_or_2_nl;
  wire[0:0] for_for_for_if_for_for_for_if_or_3_nl;
  wire[0:0] for_for_for_else_mux_5_nl;
  wire[0:0] for_for_for_else_if_for_for_for_else_if_or_1_nl;
  wire[0:0] for_for_for_else_else_mux_1_nl;
  wire[0:0] for_for_for_else_else_else_for_for_for_else_else_else_or_1_nl;
  wire[0:0] for_for_for_else_else_if_for_for_for_else_else_if_or_1_nl;
  wire[0:0] for_for_for_if_for_for_for_if_or_4_nl;
  wire[0:0] for_for_for_else_mux_7_nl;
  wire[0:0] for_for_for_else_if_for_for_for_else_if_or_nl;
  wire[0:0] for_for_for_else_else_mux_nl;
  wire[0:0] for_for_for_else_else_else_for_for_for_else_else_else_or_nl;
  wire[0:0] for_for_for_else_else_if_for_for_for_else_else_if_or_nl;
  wire[0:0] for_for_for_if_for_for_for_if_or_5_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [23:0] nl_PixelAccumulator_run_output_pxl_serial_rsci_inst_output_pxl_serial_rsci_idat;
  assign nl_PixelAccumulator_run_output_pxl_serial_rsci_inst_output_pxl_serial_rsci_idat
      = {output_pxl_serial_rsci_idat_23 , output_pxl_serial_rsci_idat_22 , output_pxl_serial_rsci_idat_21
      , output_pxl_serial_rsci_idat_20 , output_pxl_serial_rsci_idat_19 , output_pxl_serial_rsci_idat_18
      , output_pxl_serial_rsci_idat_17 , output_pxl_serial_rsci_idat_16 , output_pxl_serial_rsci_idat_15
      , output_pxl_serial_rsci_idat_14 , output_pxl_serial_rsci_idat_13 , output_pxl_serial_rsci_idat_12
      , output_pxl_serial_rsci_idat_11 , output_pxl_serial_rsci_idat_10 , output_pxl_serial_rsci_idat_9
      , output_pxl_serial_rsci_idat_8 , output_pxl_serial_rsci_idat_7 , output_pxl_serial_rsci_idat_6
      , output_pxl_serial_rsci_idat_5 , output_pxl_serial_rsci_idat_4 , output_pxl_serial_rsci_idat_3
      , output_pxl_serial_rsci_idat_2 , output_pxl_serial_rsci_idat_1 , output_pxl_serial_rsci_idat_0};
  PixelAccumulator_run_accumulator_parms_rsci PixelAccumulator_run_accumulator_parms_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .accumulator_parms_rsc_dat(accumulator_parms_rsc_dat),
      .accumulator_parms_rsc_vld(accumulator_parms_rsc_vld),
      .accumulator_parms_rsc_rdy(accumulator_parms_rsc_rdy),
      .run_wen(run_wen),
      .accumulator_parms_rsci_oswt(reg_accumulator_parms_rsci_oswt_cse),
      .accumulator_parms_rsci_wen_comp(accumulator_parms_rsci_wen_comp),
      .accumulator_parms_rsci_idat_mxwt(accumulator_parms_rsci_idat_mxwt)
    );
  PixelAccumulator_run_pxl_sample_rsci PixelAccumulator_run_pxl_sample_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .pxl_sample_rsc_dat(pxl_sample_rsc_dat),
      .pxl_sample_rsc_vld(pxl_sample_rsc_vld),
      .pxl_sample_rsc_rdy(pxl_sample_rsc_rdy),
      .run_wen(run_wen),
      .pxl_sample_rsci_oswt(reg_pxl_sample_rsci_oswt_cse),
      .pxl_sample_rsci_wen_comp(pxl_sample_rsci_wen_comp),
      .pxl_sample_rsci_idat_mxwt(pxl_sample_rsci_idat_mxwt)
    );
  PixelAccumulator_run_output_pxl_serial_rsci PixelAccumulator_run_output_pxl_serial_rsci_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy),
      .run_wen(run_wen),
      .output_pxl_serial_rsci_oswt(reg_output_pxl_serial_rsci_oswt_cse),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp),
      .output_pxl_serial_rsci_idat(nl_PixelAccumulator_run_output_pxl_serial_rsci_inst_output_pxl_serial_rsci_idat[23:0])
    );
  PixelAccumulator_run_staller PixelAccumulator_run_staller_inst (
      .run_wen(run_wen),
      .accumulator_parms_rsci_wen_comp(accumulator_parms_rsci_wen_comp),
      .pxl_sample_rsci_wen_comp(pxl_sample_rsci_wen_comp),
      .output_pxl_serial_rsci_wen_comp(output_pxl_serial_rsci_wen_comp)
    );
  assign nor_8_cse = ~((for_acc_2_tmp[11]) | operator_11_false_1_equal_1_tmp);
  assign output_pxl_serial_and_cse = run_wen & (~ or_dcpl_4);
  assign nand_3_cse = ~((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4]));
  assign nor_23_cse = ~(operator_11_false_equal_tmp | (for_for_acc_1_tmp[11]));
  assign and_27_cse = (nand_3_cse | nor_23_cse | nor_8_cse | (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1!=2'b10))
      & exitL_exit_for_sva & main_stage_0_2 & run_wen;
  assign or_20_cse = operator_11_false_equal_tmp | (for_for_acc_1_tmp[11]);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_and_cse = run_wen
      & ((~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3)
      | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1) & main_stage_0_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_and_cse
      = run_wen & ((~(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_36_cse_1
      | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3))
      | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_37_cse_1
      | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2)
      & main_stage_0_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_and_2_cse
      = run_wen & main_stage_0_2;
  assign and_69_cse = (((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
      & (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1==2'b10))
      | (~ main_stage_0_2) | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1)
      & run_wen;
  assign nor_12_nl = ~((for_for_for_samps_10_0_sva_2[10]) | ((for_for_for_samps_10_0_lpi_1_dfm_1_9_0[4:0]==5'b11111)
      & operator_33_true_equal_tmp & (operator_11_false_1_acc_sdt_sva_1[6:5]==2'b00)));
  assign mux_8_nl = MUX_s_1_2_2((nor_12_nl), (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[0]),
      lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[1]);
  assign and_81_cse = (~ (mux_8_nl)) & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_and_2_cse;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_239_tmp
      = MUX1HOT_v_2_4_2(2'b01, 2'b10, lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_3,
      lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1,
      {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_36_cse_1 ,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_37_cse_1 ,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_23_cse_1 ,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3});
  assign exitL_exit_for_sva_mx0 = MUX_s_1_2_2(exitL_exit_for_sva, exit_for_lpi_1_dfm_3_mx0w0,
      main_stage_0_2);
  assign for_mux_6_nl = MUX_s_1_2_2(operator_11_false_1_equal_1_tmp, exit_for_sva_2,
      or_tmp_7);
  assign exit_for_lpi_1_dfm_3_mx0w0 = ((for_acc_2_tmp[11]) | (for_mux_6_nl)) & exit_for_for_lpi_1_dfm_3
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign lfst_exit_for_for_lpi_1_dfm_mx0 = (~(exit_for_for_lpi_1_dfm_3 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2))
      & main_stage_0_2;
  assign operator_2_false_2_operator_2_false_2_and_mdf_sva_1 = (accumulator_parms_rsci_idat_mxwt[1:0]==2'b10);
  assign operator_2_false_1_operator_2_false_1_and_mdf_sva_1 = (accumulator_parms_rsci_idat_mxwt[1:0]==2'b01);
  assign operator_2_false_operator_2_false_nor_mdf_sva_1 = ~((accumulator_parms_rsci_idat_mxwt[1:0]!=2'b00));
  assign exit_for_for_for_lpi_1_dfm_1 = (for_for_for_samps_10_0_sva_2[10]) | exit_for_for_for_sva_1;
  assign accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0 = MUX_s_1_2_2((accumulator_parms_crt_lpi_1_dfm_12_11[0]),
      (accumulator_parms_rsci_idat_mxwt[0]), exitL_exit_for_sva);
  assign accumulator_parms_crt_lpi_1_dfm_12_11_mx2_1 = MUX_s_1_2_2((accumulator_parms_crt_lpi_1_dfm_12_11[1]),
      (accumulator_parms_rsci_idat_mxwt[1]), exitL_exit_for_sva);
  assign nl_for_for_for_samps_10_0_sva_2 = conv_u2s_10_11(for_for_for_samps_10_0_lpi_1_dfm_1_9_0)
      + 11'b00000000001;
  assign for_for_for_samps_10_0_sva_2 = nl_for_for_for_samps_10_0_sva_2[10:0];
  assign operator_33_true_equal_tmp = (for_for_for_samps_10_0_lpi_1_dfm_1_9_0[9:5])
      == (operator_11_false_1_acc_sdt_sva_1[4:0]);
  assign exit_for_for_for_sva_1 = (for_for_for_samps_10_0_lpi_1_dfm_1_9_0[4:0]==5'b11111)
      & operator_33_true_equal_tmp & (operator_11_false_1_acc_sdt_sva_1[6:5]==2'b00);
  assign nl_operator_11_false_1_acc_sdt_sva_1 = conv_u2u_6_7({mgc_qr_10_lpi_1_dfm_1_mx0
      , 1'b0 , mgc_qr_8_lpi_1_dfm_1_mx0 , 1'b0 , mgc_qr_6_lpi_1_dfm_1_mx0 , operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm_mx0})
      + 7'b1111111;
  assign operator_11_false_1_acc_sdt_sva_1 = nl_operator_11_false_1_acc_sdt_sva_1[6:0];
  assign nor_1_nl = ~(operator_2_false_2_operator_2_false_2_and_mdf_sva_1 | operator_2_false_1_operator_2_false_1_and_mdf_sva_1
      | operator_2_false_operator_2_false_nor_mdf_sva_1);
  assign mgc_qr_10_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(mgc_qr_10_lpi_1_dfm_1, (nor_1_nl),
      exitL_exit_for_sva);
  assign mgc_qr_8_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(mgc_qr_8_lpi_1_dfm_1, operator_2_false_2_operator_2_false_2_and_mdf_sva_1,
      exitL_exit_for_sva);
  assign mgc_qr_6_lpi_1_dfm_1_mx0 = MUX_s_1_2_2(mgc_qr_6_lpi_1_dfm_1, operator_2_false_1_operator_2_false_1_and_mdf_sva_1,
      exitL_exit_for_sva);
  assign operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm_mx0 = MUX_s_1_2_2(operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm,
      operator_2_false_operator_2_false_nor_mdf_sva_1, exitL_exit_for_sva);
  assign nl_for_acc_2_tmp = conv_u2s_11_12(for_fy_11_0_lpi_1_dfm_1_10_0) + 12'b000000000001;
  assign for_acc_2_tmp = nl_for_acc_2_tmp[11:0];
  assign operator_11_false_1_equal_1_tmp = (for_fy_11_0_lpi_1_dfm_1_10_0) == (operator_12_true_return_10_0_lpi_1_dfm_mx0);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_nl = ~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1;
  assign lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_3
      = MUX_v_2_2_2(2'b00, lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1,
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_nl));
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2
      = (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1==2'b10);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1
      = (~ (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_3[1]))
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign exit_for_for_lpi_1_dfm_3 = or_20_cse & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_36_cse_1
      = (~ exit_for_for_for_lpi_1_dfm_1) & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_37_cse_1
      = exit_for_for_for_lpi_1_dfm_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_23_cse_1
      = (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_3[1])
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_4
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_239_tmp
      & (signext_2_1(~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1))
      & ({{1{lfst_exit_for_for_lpi_1_dfm_mx0}}, lfst_exit_for_for_lpi_1_dfm_mx0});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3
      = (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1==2'b11);
  assign nl_operator_12_true_acc_nl = (~ (accumulator_parms_rsci_idat_mxwt[23:13]))
      + (accumulator_parms_rsci_idat_mxwt[34:24]);
  assign operator_12_true_acc_nl = nl_operator_12_true_acc_nl[10:0];
  assign operator_12_true_return_10_0_lpi_1_dfm_mx0 = MUX_v_11_2_2(operator_12_true_return_10_0_lpi_1_dfm,
      (operator_12_true_acc_nl), exitL_exit_for_sva);
  assign nl_for_for_acc_1_tmp = conv_u2s_11_12(for_for_fx_11_0_lpi_1_dfm_1_10_0)
      + 12'b000000000001;
  assign for_for_acc_1_tmp = nl_for_for_acc_1_tmp[11:0];
  assign operator_11_false_equal_tmp = (for_for_fx_11_0_lpi_1_dfm_1_10_0) == (operator_11_false_return_10_0_lpi_1_dfm_mx0);
  assign nl_operator_11_false_acc_nl = (accumulator_parms_rsci_idat_mxwt[12:2]) +
      11'b11111111111;
  assign operator_11_false_acc_nl = nl_operator_11_false_acc_nl[10:0];
  assign operator_11_false_return_10_0_lpi_1_dfm_mx0 = MUX_v_11_2_2(operator_11_false_return_10_0_lpi_1_dfm,
      (operator_11_false_acc_nl), exitL_exit_for_sva);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1
      = (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4]);
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp
      = conv_u2s_4_5(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_i_4_0_lpi_1_3_0)
      + 5'b11111;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp =
      nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4:0];
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp
      = conv_u2s_4_5(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_i_4_0_lpi_1_3_0)
      + 5'b11111;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp
      = nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4:0];
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp
      = conv_u2s_4_5(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_4_0_lpi_1_3_0)
      + 5'b11111;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp
      = nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4:0];
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_14_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_14_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_14_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_12_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_13_lpi_1;
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp
      = ({(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_14_nl)
      , (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_12_nl)
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_12_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_11_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_10_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_9_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_8_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_7_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_6_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_5_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_4_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_3_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_2_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_1_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_0_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_14_lpi_1})
      + ({1'b1 , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1) , 2'b10})
      + 17'b00000000000000001;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp
      = nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16:0];
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_14_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_14_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_14_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_12_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_13_lpi_1;
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp
      = ({(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_14_nl)
      , (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_12_nl)
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_12_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_11_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_10_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_9_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_8_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_7_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_6_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_5_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_4_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_3_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_2_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_1_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_0_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_14_lpi_1})
      + ({1'b1 , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1) , 2'b10})
      + 17'b00000000000000001;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp
      = nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16:0];
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_14_nl =
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_14_lpi_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_14_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_12_nl =
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_13_lpi_1;
  assign nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp
      = ({(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_14_nl)
      , (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_12_nl) ,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_12_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_11_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_10_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_9_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_8_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_7_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_6_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_5_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_4_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_3_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_2_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_1_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_0_sva_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_14_lpi_1})
      + ({1'b1 , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1) ,
      (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1)
      , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1) , (~
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1) , (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1)
      , 2'b10}) + 17'b00000000000000001;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp =
      nl_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16:0];
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_12_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_12_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_11_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_11_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_10_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_10_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_9_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_9_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_8_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_8_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_7_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_7_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_6_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_6_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_5_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_5_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_4_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_4_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_3_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_3_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_2_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_2_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_1_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_1_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_0_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_0_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_12_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_12_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_11_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_11_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_10_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_10_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_9_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_9_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_8_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_8_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_7_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_7_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_6_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_6_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_5_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_5_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_4_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_4_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_3_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_3_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_2_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_2_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_1_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_1_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_0_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_0_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_12_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_12_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_11_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_11_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_10_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_10_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_9_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_9_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_8_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_8_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_7_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_7_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_6_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_6_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_5_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_5_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_4_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_4_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_3_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_3_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_2_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_2_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_1_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_1_lpi_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_0_sva_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 &
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_0_lpi_1;
  assign for_for_rounded_accuracy_col_z_lpi_1_dfm_3 = MUX1HOT_v_15_4_2((for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1[19:5]),
      (for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1[17:3]), (for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1[15:1]),
      (for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1[14:0]), {(~ for_for_for_unequal_tmp_1)
      , (~ for_for_else_3_unequal_tmp_1) , for_for_asn_17 , for_for_asn_19});
  assign for_for_rounded_accuracy_col_y_lpi_1_dfm_3 = MUX1HOT_v_15_4_2((for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1[19:5]),
      (for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1[17:3]), (for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1[15:1]),
      (for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1[14:0]), {(~ for_for_for_unequal_tmp_1)
      , (~ for_for_else_3_unequal_tmp_1) , for_for_asn_17 , for_for_asn_19});
  assign for_for_rounded_accuracy_col_x_lpi_1_dfm_3 = MUX1HOT_v_15_4_2((for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1[19:5]),
      (for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1[17:3]), (for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1[15:1]),
      (for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1[14:0]), {(~ for_for_for_unequal_tmp_1)
      , (~ for_for_else_3_unequal_tmp_1) , for_for_asn_17 , for_for_asn_19});
  assign nl_for_for_for_ac_fixed_cctor_2_sva_1 = for_for_accumulation_reg_z_lpi_1_dfm_1
      + conv_u2u_27_33(pxl_sample_rsci_idat_mxwt[80:54]);
  assign for_for_for_ac_fixed_cctor_2_sva_1 = nl_for_for_for_ac_fixed_cctor_2_sva_1[32:0];
  assign nl_for_for_for_ac_fixed_cctor_1_sva_1 = for_for_accumulation_reg_y_lpi_1_dfm_1
      + conv_u2u_27_33(pxl_sample_rsci_idat_mxwt[53:27]);
  assign for_for_for_ac_fixed_cctor_1_sva_1 = nl_for_for_for_ac_fixed_cctor_1_sva_1[32:0];
  assign nl_for_for_for_ac_fixed_cctor_sva_1 = for_for_accumulation_reg_x_lpi_1_dfm_1
      + conv_u2u_27_33(pxl_sample_rsci_idat_mxwt[26:0]);
  assign for_for_for_ac_fixed_cctor_sva_1 = nl_for_for_for_ac_fixed_cctor_sva_1[32:0];
  assign for_for_else_3_unequal_tmp_1 = ~(accumulator_parms_crt_lpi_1_dfm_12_11_mx2_1
      & (~ accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0));
  assign for_for_accumulation_reg_z_lpi_1_dfm_1_32_13_1 = MUX_v_20_2_2((for_for_for_ac_fixed_cctor_2_sva_1[32:13]),
      20'b11111111111111111111, for_for_blue_of_lpi_1_dfm_7_mx0);
  assign for_for_accumulation_reg_y_lpi_1_dfm_1_32_13_1 = MUX_v_20_2_2((for_for_for_ac_fixed_cctor_1_sva_1[32:13]),
      20'b11111111111111111111, for_for_green_of_lpi_1_dfm_7_mx0);
  assign for_for_accumulation_reg_x_lpi_1_dfm_1_32_13_1 = MUX_v_20_2_2((for_for_for_ac_fixed_cctor_sva_1[32:13]),
      20'b11111111111111111111, for_for_red_of_lpi_1_dfm_7_mx0);
  assign for_for_for_unequal_tmp_1 = ~(accumulator_parms_crt_lpi_1_dfm_12_11_mx2_1
      & accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0);
  assign for_for_for_else_if_for_for_for_else_if_or_2_nl = for_for_blue_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_2_sva_1[30]);
  assign for_for_for_else_else_else_for_for_for_else_else_else_or_2_nl = for_for_blue_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_2_sva_1[27]);
  assign for_for_for_else_else_if_for_for_for_else_else_if_or_2_nl = for_for_blue_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_2_sva_1[28]);
  assign for_for_for_else_else_mux_2_nl = MUX_s_1_2_2((for_for_for_else_else_else_for_for_for_else_else_else_or_2_nl),
      (for_for_for_else_else_if_for_for_for_else_else_if_or_2_nl), accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0);
  assign for_for_for_else_mux_3_nl = MUX_s_1_2_2((for_for_for_else_if_for_for_for_else_if_or_2_nl),
      (for_for_for_else_else_mux_2_nl), for_for_else_3_unequal_tmp_1);
  assign for_for_for_if_for_for_for_if_or_3_nl = for_for_blue_of_lpi_1_dfm_1 | (for_for_for_ac_fixed_cctor_2_sva_1[32]);
  assign for_for_blue_of_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((for_for_for_else_mux_3_nl),
      (for_for_for_if_for_for_for_if_or_3_nl), and_dcpl_7);
  assign for_for_for_else_if_for_for_for_else_if_or_1_nl = for_for_green_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_1_sva_1[30]);
  assign for_for_for_else_else_else_for_for_for_else_else_else_or_1_nl = for_for_green_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_1_sva_1[27]);
  assign for_for_for_else_else_if_for_for_for_else_else_if_or_1_nl = for_for_green_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_1_sva_1[28]);
  assign for_for_for_else_else_mux_1_nl = MUX_s_1_2_2((for_for_for_else_else_else_for_for_for_else_else_else_or_1_nl),
      (for_for_for_else_else_if_for_for_for_else_else_if_or_1_nl), accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0);
  assign for_for_for_else_mux_5_nl = MUX_s_1_2_2((for_for_for_else_if_for_for_for_else_if_or_1_nl),
      (for_for_for_else_else_mux_1_nl), for_for_else_3_unequal_tmp_1);
  assign for_for_for_if_for_for_for_if_or_4_nl = for_for_green_of_lpi_1_dfm_1 | (for_for_for_ac_fixed_cctor_1_sva_1[32]);
  assign for_for_green_of_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((for_for_for_else_mux_5_nl),
      (for_for_for_if_for_for_for_if_or_4_nl), and_dcpl_7);
  assign for_for_for_else_if_for_for_for_else_if_or_nl = for_for_red_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_sva_1[30]);
  assign for_for_for_else_else_else_for_for_for_else_else_else_or_nl = for_for_red_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_sva_1[27]);
  assign for_for_for_else_else_if_for_for_for_else_else_if_or_nl = for_for_red_of_lpi_1_dfm_1
      | (for_for_for_ac_fixed_cctor_sva_1[28]);
  assign for_for_for_else_else_mux_nl = MUX_s_1_2_2((for_for_for_else_else_else_for_for_for_else_else_else_or_nl),
      (for_for_for_else_else_if_for_for_for_else_else_if_or_nl), accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0);
  assign for_for_for_else_mux_7_nl = MUX_s_1_2_2((for_for_for_else_if_for_for_for_else_if_or_nl),
      (for_for_for_else_else_mux_nl), for_for_else_3_unequal_tmp_1);
  assign for_for_for_if_for_for_for_if_or_5_nl = for_for_red_of_lpi_1_dfm_1 | (for_for_for_ac_fixed_cctor_sva_1[32]);
  assign for_for_red_of_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((for_for_for_else_mux_7_nl),
      (for_for_for_if_for_for_for_if_or_5_nl), and_dcpl_7);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_94_cse_1
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_23_cse_1
      | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3;
  assign for_for_for_and_2_tmp_1 = for_for_blue_of_lpi_1_dfm_7_mx0 & exit_for_for_for_lpi_1_dfm_1;
  assign for_for_for_and_1_tmp_1 = for_for_green_of_lpi_1_dfm_7_mx0 & exit_for_for_for_lpi_1_dfm_1;
  assign for_for_for_and_tmp_1 = for_for_red_of_lpi_1_dfm_7_mx0 & exit_for_for_for_lpi_1_dfm_1;
  assign for_for_asn_17 = accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0 & for_for_for_unequal_tmp_1;
  assign for_for_asn_19 = (~ accumulator_parms_crt_lpi_1_dfm_12_11_mx1_0) & for_for_else_3_unequal_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 = (~
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16]))
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484 = (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16])
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 = (~
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16]))
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488 = (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16])
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 = (~
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16]))
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492 = (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16])
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign for_mux_tmp = MUX_v_2_2_2(accumulator_parms_crt_lpi_1_dfm_12_11, (accumulator_parms_rsci_idat_mxwt[1:0]),
      exitL_exit_for_sva);
  assign or_tmp_7 = nor_23_cse | (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1!=2'b10)
      | (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1);
  assign or_dcpl_2 = (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1!=2'b10);
  assign or_dcpl_4 = (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1)
      | or_dcpl_2 | (~ main_stage_0_2);
  assign and_dcpl_7 = (for_mux_tmp==2'b11);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_accumulator_parms_rsci_oswt_cse <= 1'b0;
      reg_output_pxl_serial_rsci_oswt_cse <= 1'b0;
      reg_pxl_sample_rsci_oswt_cse <= 1'b0;
      lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1
          <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      for_for_blue_of_lpi_1_dfm_1 <= 1'b0;
      for_for_green_of_lpi_1_dfm_1 <= 1'b0;
      for_for_red_of_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_accumulator_parms_rsci_oswt_cse <= MUX_s_1_2_2(exitL_exit_for_sva, (nor_nl),
          main_stage_0_2);
      reg_output_pxl_serial_rsci_oswt_cse <= ~ or_dcpl_4;
      reg_pxl_sample_rsci_oswt_cse <= ~(((~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1)
          | or_dcpl_2) & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_239_tmp[1])
          & main_stage_0_2);
      lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1
          <= lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_4;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 <= ((lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_4==2'b01))
          | (~((lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_4!=2'b00)));
      main_stage_0_2 <= 1'b1;
      for_for_blue_of_lpi_1_dfm_1 <= (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_5_nl)
          & lfst_exit_for_for_lpi_1_dfm_mx0;
      for_for_green_of_lpi_1_dfm_1 <= (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_4_nl)
          & lfst_exit_for_for_lpi_1_dfm_mx0;
      for_for_red_of_lpi_1_dfm_1 <= (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_3_nl)
          & lfst_exit_for_for_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      output_pxl_serial_rsci_idat_23 <= 1'b0;
      output_pxl_serial_rsci_idat_0 <= 1'b0;
      output_pxl_serial_rsci_idat_22 <= 1'b0;
      output_pxl_serial_rsci_idat_1 <= 1'b0;
      output_pxl_serial_rsci_idat_21 <= 1'b0;
      output_pxl_serial_rsci_idat_2 <= 1'b0;
      output_pxl_serial_rsci_idat_20 <= 1'b0;
      output_pxl_serial_rsci_idat_3 <= 1'b0;
      output_pxl_serial_rsci_idat_19 <= 1'b0;
      output_pxl_serial_rsci_idat_4 <= 1'b0;
      output_pxl_serial_rsci_idat_18 <= 1'b0;
      output_pxl_serial_rsci_idat_5 <= 1'b0;
      output_pxl_serial_rsci_idat_17 <= 1'b0;
      output_pxl_serial_rsci_idat_6 <= 1'b0;
      output_pxl_serial_rsci_idat_16 <= 1'b0;
      output_pxl_serial_rsci_idat_7 <= 1'b0;
      output_pxl_serial_rsci_idat_15 <= 1'b0;
      output_pxl_serial_rsci_idat_8 <= 1'b0;
      output_pxl_serial_rsci_idat_14 <= 1'b0;
      output_pxl_serial_rsci_idat_9 <= 1'b0;
      output_pxl_serial_rsci_idat_13 <= 1'b0;
      output_pxl_serial_rsci_idat_10 <= 1'b0;
      output_pxl_serial_rsci_idat_12 <= 1'b0;
      output_pxl_serial_rsci_idat_11 <= 1'b0;
    end
    else if ( output_pxl_serial_and_cse ) begin
      output_pxl_serial_rsci_idat_23 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_0 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_22 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_1 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_21 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_2 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_20 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_3 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_19 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_4 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_18 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_5 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_17 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_6 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_16 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1;
      output_pxl_serial_rsci_idat_7 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1;
      output_pxl_serial_rsci_idat_15 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_8 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_14 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_9 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_13 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_10 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_12 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
      output_pxl_serial_rsci_idat_11 <= ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exit_for_sva <= 1'b1;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 <= 1'b0;
    end
    else if ( ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_and_2_cse
        ) begin
      exitL_exit_for_sva <= exitL_exit_for_sva_mx0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1 <=
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_65_nl)
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1 <=
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_64_nl)
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 <= (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_63_nl)
          | ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumulator_parms_crt_lpi_1_dfm_12_11 <= 2'b00;
    end
    else if ( run_wen & (~(((for_acc_2_tmp[11]) | operator_11_false_1_equal_1_tmp)
        & (~(nor_23_cse | (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1!=2'b10)
        | nand_3_cse)))) & main_stage_0_2 & exitL_exit_for_sva ) begin
      accumulator_parms_crt_lpi_1_dfm_12_11 <= accumulator_parms_rsci_idat_mxwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_for_samps_10_0_lpi_1_dfm_1_9_0 <= 10'b0000000000;
    end
    else if ( (~((mux_nl) & main_stage_0_2)) & run_wen ) begin
      for_for_for_samps_10_0_lpi_1_dfm_1_9_0 <= MUX_v_10_2_2(10'b0000000000, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_96_nl),
          lfst_exit_for_for_lpi_1_dfm_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_for_for_for_sva <= 1'b0;
    end
    else if ( run_wen & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_239_tmp[1])
        & main_stage_0_2 & (~ (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[1]))
        ) begin
      exit_for_for_for_sva <= exit_for_for_for_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      mgc_qr_10_lpi_1_dfm_1 <= 1'b0;
      mgc_qr_8_lpi_1_dfm_1 <= 1'b0;
      mgc_qr_6_lpi_1_dfm_1 <= 1'b0;
      operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm <= 1'b0;
      operator_12_true_return_10_0_lpi_1_dfm <= 11'b00000000000;
      operator_11_false_return_10_0_lpi_1_dfm <= 11'b00000000000;
    end
    else if ( and_27_cse ) begin
      mgc_qr_10_lpi_1_dfm_1 <= mgc_qr_10_lpi_1_dfm_1_mx0;
      mgc_qr_8_lpi_1_dfm_1 <= mgc_qr_8_lpi_1_dfm_1_mx0;
      mgc_qr_6_lpi_1_dfm_1 <= mgc_qr_6_lpi_1_dfm_1_mx0;
      operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm <= operator_2_false_operator_2_false_nor_mdf_lpi_1_dfm_mx0;
      operator_12_true_return_10_0_lpi_1_dfm <= operator_12_true_return_10_0_lpi_1_dfm_mx0;
      operator_11_false_return_10_0_lpi_1_dfm <= operator_11_false_return_10_0_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exit_for_sva_2 <= 1'b0;
    end
    else if ( run_wen & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
        & (~ (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[0]))
        & or_20_cse & (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[1])
        & main_stage_0_2 ) begin
      exit_for_sva_2 <= operator_11_false_1_equal_1_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_fy_11_0_lpi_1_dfm_1_10_0 <= 11'b00000000000;
    end
    else if ( (((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
        & (~ (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[0]))
        & or_20_cse & (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[1]))
        | (exitL_exit_for_sva & (~ main_stage_0_2))) & run_wen ) begin
      for_fy_11_0_lpi_1_dfm_1_10_0 <= MUX_v_11_2_2(11'b00000000000, (for_acc_2_tmp[10:0]),
          (for_not_20_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_fx_11_0_lpi_1_dfm_1_10_0 <= 11'b00000000000;
    end
    else if ( (~((~((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
        & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
        & (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1==2'b10)))
        & main_stage_0_2)) & run_wen ) begin
      for_for_fx_11_0_lpi_1_dfm_1_10_0 <= MUX_v_11_2_2(11'b00000000000, (for_for_for_for_for_for_mux_nl),
          (for_for_for_for_not_nl));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_14_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_7_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_14_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_7_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_14_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_13_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_0_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_1_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_12_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_2_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 <=
          1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_11_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_3_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_10_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_4_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_9_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_5_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_8_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_6_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_7_lpi_1 <= 1'b0;
    end
    else if ( ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_and_cse
        ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_77_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_76_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_24_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_16_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_78_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_23_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_79_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_22_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_80_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_21_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_81_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_20_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_82_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_19_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_83_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_18_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_84_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_17_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_47_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_46_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_54_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_48_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_53_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_49_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_52_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_50_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_51_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_85_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_55_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_25_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_86_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_56_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_26_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_87_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_57_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_27_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_88_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_58_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_28_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_89_nl),
          (~ (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16])),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_59_nl),
          (~ (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16])),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_29_nl),
          (~ (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16])),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_14_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_106_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_14_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_61_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_14_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_12_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_107_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_13_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_62_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_12_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_11_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_60_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_13_12_lpi_1[1]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_75_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_2_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_74_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_3_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_12_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_63_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_10_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_10_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_112_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_2_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_73_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_9_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_0_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_108_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_11_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_64_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_8_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_9_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_3_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_72_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_7_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_1_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_10_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_65_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_6_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_8_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_111_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_4_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_71_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_5_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_2_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_109_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_9_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_66_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_4_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_7_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_5_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_70_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_3_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_3_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_8_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_67_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_2_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_6_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_110_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_6_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_69_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_1_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_4_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_7_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_68_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_and_psp_5_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_482 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_484});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_14_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_98_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_14_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_31_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_14_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_12_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_99_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_13_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_32_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_12_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_11_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_30_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_13_12_lpi_1[1]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_45_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_2_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_44_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_3_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_12_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_33_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_10_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_10_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_104_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_2_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_43_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_9_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_0_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_100_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_11_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_34_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_8_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_9_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_3_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_42_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_7_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_1_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_10_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_35_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_6_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_8_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_103_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_4_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_41_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_5_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_2_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_101_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_9_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_36_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_4_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_7_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_5_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_40_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_3_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_3_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_8_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_37_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_2_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_6_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_102_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_6_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_39_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_1_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_4_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_7_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_38_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_and_psp_5_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_486 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_488});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_14_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_90_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_14_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_1_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_14_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_12_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_91_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_13_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_2_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_12_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_11_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_13_12_lpi_1[1]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_0_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_15_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_2_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_1_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_14_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_3_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_12_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_3_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_10_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_10_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_96_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_2_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_13_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_9_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_0_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 <=
          MUX_s_1_2_2((for_for_for_for_for_for_and_92_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_11_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_4_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_8_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_9_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_3_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_12_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_7_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_1_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_10_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_5_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_6_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_8_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_95_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_4_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_11_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_5_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_2_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_93_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_9_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_6_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_4_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_7_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_5_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_10_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_3_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_3_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_8_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_7_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_2_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_6_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 <= MUX_s_1_2_2((for_for_for_for_for_for_and_94_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_6_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_9_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_1_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_4_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_7_lpi_1 <= MUX1HOT_s_1_3_2((for_for_for_for_for_for_and_8_nl),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_nl),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_psp_5_sva_1,
          {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1 ,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_490 , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_asn_492});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_4_0_lpi_1_3_0
          <= 4'b0000;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_i_4_0_lpi_1_3_0
          <= 4'b0000;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_i_4_0_lpi_1_3_0
          <= 4'b0000;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_14_lpi_1 <= 1'b0;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_13_12_lpi_1 <=
          2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_13_12_lpi_1 <=
          2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_13_12_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_11_10_lpi_1 <=
          2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_11_10_lpi_1 <=
          2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_11_10_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_9_8_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_9_8_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_9_8_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_7_6_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_7_6_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_7_6_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_5_4_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_5_4_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_5_4_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_3_2_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_3_2_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_3_2_lpi_1 <= 2'b00;
    end
    else if ( ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_and_cse
        ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_i_4_0_lpi_1_3_0
          <= MUX_v_4_2_2(4'b1110, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[3:0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_i_4_0_lpi_1_3_0
          <= MUX_v_4_2_2(4'b1110, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[3:0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_i_4_0_lpi_1_3_0
          <= MUX_v_4_2_2(4'b1110, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[3:0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_14_lpi_1 <= MUX_s_1_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[14]),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_13_12_lpi_1[0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_14_lpi_1 <= MUX_s_1_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[14]),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_13_12_lpi_1[0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_14_lpi_1 <= MUX_s_1_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[14]),
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_13_12_lpi_1[0]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_13_12_lpi_1 <=
          MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[13:12]), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_11_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_13_12_lpi_1 <=
          MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[13:12]), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_11_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_13_12_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[13:12]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_11_10_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_11_10_lpi_1 <=
          MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[11:10]), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_9_8_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_11_10_lpi_1 <=
          MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[11:10]), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_9_8_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_11_10_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[11:10]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_9_8_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_9_8_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[9:8]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_7_6_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_9_8_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[9:8]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_7_6_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_9_8_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[9:8]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_7_6_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_7_6_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[7:6]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_5_4_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_7_6_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[7:6]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_5_4_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_7_6_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[7:6]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_5_4_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_5_4_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[5:4]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_3_2_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_5_4_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[5:4]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_3_2_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_5_4_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[5:4]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_3_2_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_3_2_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_z_lpi_1_dfm_3[3:2]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_1_0_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_3_2_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_y_lpi_1_dfm_3[3:2]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_1_0_lpi_1,
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_3_2_lpi_1 <= MUX_v_2_2_2((for_for_rounded_accuracy_col_x_lpi_1_dfm_3[3:2]),
          ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_1_0_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      for_for_accumulation_reg_z_lpi_1_dfm_1 <= 33'b000000000000000000000000000000000;
      for_for_accumulation_reg_y_lpi_1_dfm_1 <= 33'b000000000000000000000000000000000;
      for_for_accumulation_reg_x_lpi_1_dfm_1 <= 33'b000000000000000000000000000000000;
    end
    else if ( and_69_cse ) begin
      for_for_accumulation_reg_z_lpi_1_dfm_1 <= MUX_v_33_2_2(33'b000000000000000000000000000000000,
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_2_nl),
          lfst_exit_for_for_lpi_1_dfm_mx0);
      for_for_accumulation_reg_y_lpi_1_dfm_1 <= MUX_v_33_2_2(33'b000000000000000000000000000000000,
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_1_nl),
          lfst_exit_for_for_lpi_1_dfm_mx0);
      for_for_accumulation_reg_x_lpi_1_dfm_1 <= MUX_v_33_2_2(33'b000000000000000000000000000000000,
          (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_nl),
          lfst_exit_for_for_lpi_1_dfm_mx0);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_1_0_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_1_0_lpi_1 <= 2'b00;
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_1_0_lpi_1 <= 2'b00;
    end
    else if ( and_81_cse ) begin
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_1_0_lpi_1 <= MUX_v_2_2_2(2'b00,
          (for_for_rounded_accuracy_col_z_lpi_1_dfm_3[1:0]), (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_174_nl));
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_1_0_lpi_1 <= MUX_v_2_2_2(2'b00,
          (for_for_rounded_accuracy_col_y_lpi_1_dfm_3[1:0]), (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_175_nl));
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_1_0_lpi_1 <= MUX_v_2_2_2(2'b00,
          (for_for_rounded_accuracy_col_x_lpi_1_dfm_3[1:0]), (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_37_nl));
    end
  end
  assign nor_nl = ~(nor_8_cse | or_tmp_7);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_10_nl
      = for_for_blue_of_lpi_1_dfm_1 & exit_for_for_lpi_1_dfm_3;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_5_nl =
      MUX1HOT_s_1_3_2(for_for_blue_of_lpi_1_dfm_7_mx0, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_10_nl),
      for_for_blue_of_lpi_1_dfm_1, {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_94_cse_1});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_9_nl
      = for_for_green_of_lpi_1_dfm_1 & exit_for_for_lpi_1_dfm_3;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_4_nl =
      MUX1HOT_s_1_3_2(for_for_green_of_lpi_1_dfm_7_mx0, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_9_nl),
      for_for_green_of_lpi_1_dfm_1, {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_94_cse_1});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_8_nl
      = for_for_red_of_lpi_1_dfm_1 & exit_for_for_lpi_1_dfm_3;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_3_nl =
      MUX1HOT_s_1_3_2(for_for_red_of_lpi_1_dfm_7_mx0, (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_8_nl),
      for_for_red_of_lpi_1_dfm_1, {ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_94_cse_1});
  assign for_for_for_for_for_for_and_113_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_65_nl =
      MUX_s_1_2_2((for_for_for_for_for_for_and_113_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3);
  assign for_for_for_for_for_for_and_105_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_64_nl =
      MUX_s_1_2_2((for_for_for_for_for_for_and_105_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3);
  assign for_for_for_for_for_for_and_97_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_63_nl =
      MUX_s_1_2_2((for_for_for_for_for_for_and_97_nl), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_3);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux_96_nl
      = MUX_v_10_2_2((for_for_for_samps_10_0_sva_2[9:0]), ({{9{exit_for_for_lpi_1_dfm_3}},
      exit_for_for_lpi_1_dfm_3}), ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1);
  assign nand_14_nl = ~((~((for_for_for_samps_10_0_lpi_1_dfm_1_9_0[4:0]==5'b11111)
      & operator_33_true_equal_tmp & (operator_11_false_1_acc_sdt_sva_1[6:5]==2'b00)))
      & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1);
  assign and_89_nl = (~((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_acc_1_tmp[4])
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_acc_1_tmp[4])
      & (~ (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[0]))))
      & (exit_for_for_for_sva | (~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1));
  assign mux_nl = MUX_s_1_2_2((nand_14_nl), (and_89_nl), lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1[1]);
  assign for_not_20_nl = ~ exitL_exit_for_sva_mx0;
  assign for_for_and_9_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_16_svs_1
      & (lfst_exit_ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_lpi_1_dfm_1==2'b10)
      & lfst_exit_for_for_lpi_1_dfm_mx0;
  assign for_for_for_for_for_for_mux_nl = MUX_v_11_2_2(({{10{exit_for_lpi_1_dfm_3_mx0w0}},
      exit_for_lpi_1_dfm_3_mx0w0}), (for_for_acc_1_tmp[10:0]), for_for_and_9_nl);
  assign for_for_for_for_not_nl = ~ exitL_exit_for_sva_mx0;
  assign for_for_for_for_for_for_and_77_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_76_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_24_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_16_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_78_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_23_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_79_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_22_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_80_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_21_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_81_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_20_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_82_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_19_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_83_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_18_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_84_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_17_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_47_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_46_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_54_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_48_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_53_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_49_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_52_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_50_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_51_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_85_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_55_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_25_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_86_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_56_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_26_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_87_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_57_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_27_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_88_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_58_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_28_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_89_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_r_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_59_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_r_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_29_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_r_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_106_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_61_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_14_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[14]);
  assign for_for_for_for_for_for_and_107_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_62_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_12_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[13]);
  assign for_for_for_for_for_for_and_60_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_75_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_2_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[0]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_14_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_74_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_mux_3_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[1]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_z_15_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_63_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_10_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[12]);
  assign for_for_for_for_for_for_and_112_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_73_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_9_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[2]);
  assign for_for_for_for_for_for_and_108_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_64_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_8_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[11]);
  assign for_for_for_for_for_for_and_72_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_7_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_0_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[3]);
  assign for_for_for_for_for_for_and_65_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_6_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[10]);
  assign for_for_for_for_for_for_and_111_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_71_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_5_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[4]);
  assign for_for_for_for_for_for_and_109_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_66_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_4_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[9]);
  assign for_for_for_for_for_for_and_70_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_3_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_2_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[5]);
  assign for_for_for_for_for_for_and_67_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_2_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[8]);
  assign for_for_for_for_for_for_and_110_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_69_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_1_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[6]);
  assign for_for_for_for_for_for_and_68_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_d_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_if_and_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_mask_d_4_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_2_for_t_acc_tmp[7]);
  assign for_for_for_for_for_for_and_98_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_31_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_14_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[14]);
  assign for_for_for_for_for_for_and_99_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_32_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_12_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[13]);
  assign for_for_for_for_for_for_and_30_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_45_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_2_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[0]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_14_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_44_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_mux_3_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[1]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_z_15_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_33_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_10_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[12]);
  assign for_for_for_for_for_for_and_104_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_43_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_9_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[2]);
  assign for_for_for_for_for_for_and_100_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_34_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_8_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[11]);
  assign for_for_for_for_for_for_and_42_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_7_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_0_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[3]);
  assign for_for_for_for_for_for_and_35_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_6_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[10]);
  assign for_for_for_for_for_for_and_103_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_41_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_5_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[4]);
  assign for_for_for_for_for_for_and_101_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_36_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_4_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[9]);
  assign for_for_for_for_for_for_and_40_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_3_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_2_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[5]);
  assign for_for_for_for_for_for_and_37_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_2_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[8]);
  assign for_for_for_for_for_for_and_102_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_39_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_1_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[6]);
  assign for_for_for_for_for_for_and_38_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_d_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_if_and_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_mask_d_4_lpi_1
      & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_1_for_t_acc_tmp[7]);
  assign for_for_for_for_for_for_and_90_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_1_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_14_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_14_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[14]);
  assign for_for_for_for_for_for_and_91_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_2_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_13_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_12_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[13]);
  assign for_for_for_for_for_for_and_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_15_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_0_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_2_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[0]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_14_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_14_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_1_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_mux_3_nl = MUX_s_1_2_2((ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[1]),
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_z_15_lpi_1, ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[16]);
  assign for_for_for_for_for_for_and_3_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_12_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_10_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[12]);
  assign for_for_for_for_for_for_and_96_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_13_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_2_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_9_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[2]);
  assign for_for_for_for_for_for_and_92_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_4_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_11_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_8_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[11]);
  assign for_for_for_for_for_for_and_12_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_3_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_7_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_0_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[3]);
  assign for_for_for_for_for_for_and_5_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_10_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_6_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[10]);
  assign for_for_for_for_for_for_and_95_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_11_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_4_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_5_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[4]);
  assign for_for_for_for_for_for_and_93_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_6_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_9_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_4_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[9]);
  assign for_for_for_for_for_for_and_10_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_5_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_3_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_2_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[5]);
  assign for_for_for_for_for_for_and_7_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_8_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_2_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[8]);
  assign for_for_for_for_for_for_and_94_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign for_for_for_for_for_for_and_9_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_6_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_1_nl
      = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 &
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[6]);
  assign for_for_for_for_for_for_and_8_nl = ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_d_7_lpi_1
      & (~ exit_for_for_for_lpi_1_dfm_1);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_if_and_nl =
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_mask_d_4_lpi_1 & (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_t_acc_tmp[7]);
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_172_nl =
      (~ for_for_for_and_2_tmp_1) & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_173_nl =
      for_for_for_and_2_tmp_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_2_nl =
      MUX1HOT_v_33_3_2(for_for_for_ac_fixed_cctor_2_sva_1, 33'b111111111111111111111111111111110,
      ({{32{exit_for_for_lpi_1_dfm_3}}, exit_for_for_lpi_1_dfm_3}), {(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_172_nl)
      , (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_173_nl)
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_170_nl =
      (~ for_for_for_and_1_tmp_1) & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_171_nl =
      for_for_for_and_1_tmp_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_1_nl =
      MUX1HOT_v_33_3_2(for_for_for_ac_fixed_cctor_1_sva_1, 33'b111111111111111111111111111111110,
      ({{32{exit_for_for_lpi_1_dfm_3}}, exit_for_for_lpi_1_dfm_3}), {(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_170_nl)
      , (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_171_nl)
      , ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_168_nl =
      (~ for_for_for_and_tmp_1) & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_169_nl =
      for_for_for_and_tmp_1 & ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_or_tmp_1;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_mux1h_nl = MUX1HOT_v_33_3_2(for_for_for_ac_fixed_cctor_sva_1,
      33'b111111111111111111111111111111110, ({{32{exit_for_for_lpi_1_dfm_3}}, exit_for_for_lpi_1_dfm_3}),
      {(ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_168_nl) ,
      (ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_169_nl) ,
      ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_and_22_cse_1});
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_174_nl =
      ~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_175_nl =
      ~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;
  assign ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_not_37_nl =
      ~ ac_math_ac_sqrt_15_1_AC_TRN_AC_WRAP_15_1_AC_TRN_AC_WRAP_for_equal_tmp_2;

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [14:0] MUX1HOT_v_15_4_2;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [3:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    MUX1HOT_v_15_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [32:0] MUX1HOT_v_33_3_2;
    input [32:0] input_2;
    input [32:0] input_1;
    input [32:0] input_0;
    input [2:0] sel;
    reg [32:0] result;
  begin
    result = input_0 & {33{sel[0]}};
    result = result | ( input_1 & {33{sel[1]}});
    result = result | ( input_2 & {33{sel[2]}});
    MUX1HOT_v_33_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [32:0] MUX_v_33_2_2;
    input [32:0] input_0;
    input [32:0] input_1;
    input [0:0] sel;
    reg [32:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_33_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2s_11_12 =  {1'b0, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_27_33 ;
    input [26:0]  vector ;
  begin
    conv_u2u_27_33 = {{6{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ParamsDeserializer
// ------------------------------------------------------------------


module ParamsDeserializer (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      qbuffer_params_rsc_dat, qbuffer_params_rsc_vld, qbuffer_params_rsc_rdy, render_params_rsc_dat,
      render_params_rsc_vld, render_params_rsc_rdy, accum_params_rsc_dat, accum_params_rsc_vld,
      accum_params_rsc_rdy, quad_serial_out_rsc_dat, quad_serial_out_rsc_vld, quad_serial_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [11:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [56:0] qbuffer_params_rsc_dat;
  output qbuffer_params_rsc_vld;
  input qbuffer_params_rsc_rdy;
  output [419:0] render_params_rsc_dat;
  output render_params_rsc_vld;
  input render_params_rsc_rdy;
  output [419:0] accum_params_rsc_dat;
  output accum_params_rsc_vld;
  input accum_params_rsc_rdy;
  output [376:0] quad_serial_out_rsc_dat;
  output quad_serial_out_rsc_vld;
  input quad_serial_out_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ParamsDeserializer_run ParamsDeserializer_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .qbuffer_params_rsc_dat(qbuffer_params_rsc_dat),
      .qbuffer_params_rsc_vld(qbuffer_params_rsc_vld),
      .qbuffer_params_rsc_rdy(qbuffer_params_rsc_rdy),
      .render_params_rsc_dat(render_params_rsc_dat),
      .render_params_rsc_vld(render_params_rsc_vld),
      .render_params_rsc_rdy(render_params_rsc_rdy),
      .accum_params_rsc_dat(accum_params_rsc_dat),
      .accum_params_rsc_vld(accum_params_rsc_vld),
      .accum_params_rsc_rdy(accum_params_rsc_rdy),
      .quad_serial_out_rsc_dat(quad_serial_out_rsc_dat),
      .quad_serial_out_rsc_vld(quad_serial_out_rsc_vld),
      .quad_serial_out_rsc_rdy(quad_serial_out_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    QuadBuffer_64
// ------------------------------------------------------------------


module QuadBuffer_64 (
  clk, arst_n, quads_in_rsc_dat, quads_in_rsc_vld, quads_in_rsc_rdy, paramsIn_rsc_dat,
      paramsIn_rsc_vld, paramsIn_rsc_rdy, quads_out_rsc_dat, quads_out_rsc_vld, quads_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [376:0] quads_in_rsc_dat;
  input quads_in_rsc_vld;
  output quads_in_rsc_rdy;
  input [56:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [376:0] quads_out_rsc_dat;
  output quads_out_rsc_vld;
  input quads_out_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  QuadBuffer_64_run QuadBuffer_64_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsc_dat(quads_in_rsc_dat),
      .quads_in_rsc_vld(quads_in_rsc_vld),
      .quads_in_rsc_rdy(quads_in_rsc_rdy),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .quads_out_rsc_dat(quads_out_rsc_dat),
      .quads_out_rsc_vld(quads_out_rsc_vld),
      .quads_out_rsc_rdy(quads_out_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RenderLooper
// ------------------------------------------------------------------


module RenderLooper (
  clk, arst_n, render_params_rsc_dat, render_params_rsc_vld, render_params_rsc_rdy,
      render_params_out_rsc_dat, render_params_out_rsc_vld, render_params_out_rsc_rdy,
      loopIndicesOut_rsc_dat, loopIndicesOut_rsc_vld, loopIndicesOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [419:0] render_params_rsc_dat;
  input render_params_rsc_vld;
  output render_params_rsc_rdy;
  output [419:0] render_params_out_rsc_dat;
  output render_params_out_rsc_vld;
  input render_params_out_rsc_rdy;
  output [22:0] loopIndicesOut_rsc_dat;
  output loopIndicesOut_rsc_vld;
  input loopIndicesOut_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  RenderLooper_run RenderLooper_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsc_dat(render_params_rsc_dat),
      .render_params_rsc_vld(render_params_rsc_vld),
      .render_params_rsc_rdy(render_params_rsc_rdy),
      .render_params_out_rsc_dat(render_params_out_rsc_dat),
      .render_params_out_rsc_vld(render_params_out_rsc_vld),
      .render_params_out_rsc_rdy(render_params_out_rsc_rdy),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayGeneration
// ------------------------------------------------------------------


module RayGeneration (
  clk, arst_n, loopIndicesIn_rsc_dat, loopIndicesIn_rsc_vld, loopIndicesIn_rsc_rdy,
      paramsIn_rsc_dat, paramsIn_rsc_vld, paramsIn_rsc_rdy, paramsOut_rsc_dat, paramsOut_rsc_vld,
      paramsOut_rsc_rdy, rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [22:0] loopIndicesIn_rsc_dat;
  input loopIndicesIn_rsc_vld;
  output loopIndicesIn_rsc_rdy;
  input [419:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;


  // Interconnect Declarations
  wire [24:0] psq_vecMul1_run_mul_cmp_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_b;
  wire [24:0] psq_vecMul1_run_mul_cmp_1_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_1_b;
  wire [24:0] psq_vecMul1_run_mul_cmp_2_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_2_b;
  wire [24:0] psq_vecMul1_run_mul_cmp_3_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_3_b;
  wire [24:0] psq_vecMul1_run_mul_cmp_4_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_4_b;
  wire [24:0] psq_vecMul1_run_mul_cmp_5_a;
  wire [31:0] psq_vecMul1_run_mul_cmp_5_b;


  // Interconnect Declarations for Component Instantiations 
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_a)
      * $signed(psq_vecMul1_run_mul_cmp_b));
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_1_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_1_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_1_a)
      * $signed(psq_vecMul1_run_mul_cmp_1_b));
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_2_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_2_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_2_a)
      * $signed(psq_vecMul1_run_mul_cmp_2_b));
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_3_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_3_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_3_a)
      * $signed(psq_vecMul1_run_mul_cmp_3_b));
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_4_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_4_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_4_a)
      * $signed(psq_vecMul1_run_mul_cmp_4_b));
  wire [56:0] nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_5_z;
  assign nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_5_z = conv_u2u_57_57($signed(psq_vecMul1_run_mul_cmp_5_a)
      * $signed(psq_vecMul1_run_mul_cmp_5_b));
  RayGeneration_run RayGeneration_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .rayOut_rsc_dat(rayOut_rsc_dat),
      .rayOut_rsc_vld(rayOut_rsc_vld),
      .rayOut_rsc_rdy(rayOut_rsc_rdy),
      .psq_vecMul1_run_mul_cmp_a(psq_vecMul1_run_mul_cmp_a),
      .psq_vecMul1_run_mul_cmp_b(psq_vecMul1_run_mul_cmp_b),
      .psq_vecMul1_run_mul_cmp_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_z[56:0]),
      .psq_vecMul1_run_mul_cmp_1_a(psq_vecMul1_run_mul_cmp_1_a),
      .psq_vecMul1_run_mul_cmp_1_b(psq_vecMul1_run_mul_cmp_1_b),
      .psq_vecMul1_run_mul_cmp_1_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_1_z[56:0]),
      .psq_vecMul1_run_mul_cmp_2_a(psq_vecMul1_run_mul_cmp_2_a),
      .psq_vecMul1_run_mul_cmp_2_b(psq_vecMul1_run_mul_cmp_2_b),
      .psq_vecMul1_run_mul_cmp_2_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_2_z[56:0]),
      .psq_vecMul1_run_mul_cmp_3_a(psq_vecMul1_run_mul_cmp_3_a),
      .psq_vecMul1_run_mul_cmp_3_b(psq_vecMul1_run_mul_cmp_3_b),
      .psq_vecMul1_run_mul_cmp_3_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_3_z[56:0]),
      .psq_vecMul1_run_mul_cmp_4_a(psq_vecMul1_run_mul_cmp_4_a),
      .psq_vecMul1_run_mul_cmp_4_b(psq_vecMul1_run_mul_cmp_4_b),
      .psq_vecMul1_run_mul_cmp_4_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_4_z[56:0]),
      .psq_vecMul1_run_mul_cmp_5_a(psq_vecMul1_run_mul_cmp_5_a),
      .psq_vecMul1_run_mul_cmp_5_b(psq_vecMul1_run_mul_cmp_5_b),
      .psq_vecMul1_run_mul_cmp_5_z(nl_RayGeneration_run_inst_psq_vecMul1_run_mul_cmp_5_z[56:0])
    );

  function automatic [56:0] conv_u2u_57_57 ;
    input [56:0]  vector ;
  begin
    conv_u2u_57_57 = vector;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    LoopDistrib
// ------------------------------------------------------------------


module LoopDistrib (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy,
      attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld, accumalated_color_chan_in_rsc_rdy,
      attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      ray_out_loopone_rsc_dat, ray_out_loopone_rsc_vld, ray_out_loopone_rsc_rdy,
      ray_out_looptwo_rsc_dat, ray_out_looptwo_rsc_vld, ray_out_looptwo_rsc_rdy,
      ray_out_worldhit_rsc_dat, ray_out_worldhit_rsc_vld, ray_out_worldhit_rsc_rdy,
      quad_out_loopone_rsc_dat, quad_out_loopone_rsc_vld, quad_out_loopone_rsc_rdy,
      quad_out_looptwo_rsc_dat, quad_out_looptwo_rsc_vld, quad_out_looptwo_rsc_rdy,
      quad_max_outone_rsc_dat, quad_max_outone_rsc_vld, quad_max_outone_rsc_rdy,
      quad_max_outtwo_rsc_dat, quad_max_outtwo_rsc_vld, quad_max_outtwo_rsc_rdy,
      params_out_rsc_dat, params_out_rsc_vld, params_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [165:0] ray_out_loopone_rsc_dat;
  output ray_out_loopone_rsc_vld;
  input ray_out_loopone_rsc_rdy;
  output [165:0] ray_out_looptwo_rsc_dat;
  output ray_out_looptwo_rsc_vld;
  input ray_out_looptwo_rsc_rdy;
  output [165:0] ray_out_worldhit_rsc_dat;
  output ray_out_worldhit_rsc_vld;
  input ray_out_worldhit_rsc_rdy;
  output [376:0] quad_out_loopone_rsc_dat;
  output quad_out_loopone_rsc_vld;
  input quad_out_loopone_rsc_rdy;
  output [376:0] quad_out_looptwo_rsc_dat;
  output quad_out_looptwo_rsc_vld;
  input quad_out_looptwo_rsc_rdy;
  output [10:0] quad_max_outone_rsc_dat;
  output quad_max_outone_rsc_vld;
  input quad_max_outone_rsc_rdy;
  output [10:0] quad_max_outtwo_rsc_dat;
  output quad_max_outtwo_rsc_vld;
  input quad_max_outtwo_rsc_rdy;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  LoopDistrib_run LoopDistrib_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .quads_rsc_dat(quads_rsc_dat),
      .quads_rsc_vld(quads_rsc_vld),
      .quads_rsc_rdy(quads_rsc_rdy),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .ray_out_loopone_rsc_dat(ray_out_loopone_rsc_dat),
      .ray_out_loopone_rsc_vld(ray_out_loopone_rsc_vld),
      .ray_out_loopone_rsc_rdy(ray_out_loopone_rsc_rdy),
      .ray_out_looptwo_rsc_dat(ray_out_looptwo_rsc_dat),
      .ray_out_looptwo_rsc_vld(ray_out_looptwo_rsc_vld),
      .ray_out_looptwo_rsc_rdy(ray_out_looptwo_rsc_rdy),
      .ray_out_worldhit_rsc_dat(ray_out_worldhit_rsc_dat),
      .ray_out_worldhit_rsc_vld(ray_out_worldhit_rsc_vld),
      .ray_out_worldhit_rsc_rdy(ray_out_worldhit_rsc_rdy),
      .quad_out_loopone_rsc_dat(quad_out_loopone_rsc_dat),
      .quad_out_loopone_rsc_vld(quad_out_loopone_rsc_vld),
      .quad_out_loopone_rsc_rdy(quad_out_loopone_rsc_rdy),
      .quad_out_looptwo_rsc_dat(quad_out_looptwo_rsc_dat),
      .quad_out_looptwo_rsc_vld(quad_out_looptwo_rsc_vld),
      .quad_out_looptwo_rsc_rdy(quad_out_looptwo_rsc_rdy),
      .quad_max_outone_rsc_dat(quad_max_outone_rsc_dat),
      .quad_max_outone_rsc_vld(quad_max_outone_rsc_vld),
      .quad_max_outone_rsc_rdy(quad_max_outone_rsc_rdy),
      .quad_max_outtwo_rsc_dat(quad_max_outtwo_rsc_dat),
      .quad_max_outtwo_rsc_vld(quad_max_outtwo_rsc_vld),
      .quad_max_outtwo_rsc_rdy(quad_max_outtwo_rsc_rdy),
      .params_out_rsc_dat(params_out_rsc_dat),
      .params_out_rsc_vld(params_out_rsc_vld),
      .params_out_rsc_rdy(params_out_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    IntersecLoop
// ------------------------------------------------------------------


module IntersecLoop (
  clk, arst_n, quads_rsc_dat, quads_rsc_vld, quads_rsc_rdy, ray_temp_in_rsc_dat,
      ray_temp_in_rsc_vld, ray_temp_in_rsc_rdy, quad_max_in_rsc_dat, quad_max_in_rsc_vld,
      quad_max_in_rsc_rdy, quad_hit_anything_out_rsc_dat, quad_hit_anything_out_rsc_vld,
      quad_hit_anything_out_rsc_rdy, rec_quad_out_rsc_dat, rec_quad_out_rsc_vld,
      rec_quad_out_rsc_rdy, closest_so_far_out_rsc_dat, closest_so_far_out_rsc_vld,
      closest_so_far_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [376:0] quads_rsc_dat;
  input quads_rsc_vld;
  output quads_rsc_rdy;
  input [165:0] ray_temp_in_rsc_dat;
  input ray_temp_in_rsc_vld;
  output ray_temp_in_rsc_rdy;
  input [10:0] quad_max_in_rsc_dat;
  input quad_max_in_rsc_vld;
  output quad_max_in_rsc_rdy;
  output quad_hit_anything_out_rsc_dat;
  output quad_hit_anything_out_rsc_vld;
  input quad_hit_anything_out_rsc_rdy;
  output [225:0] rec_quad_out_rsc_dat;
  output rec_quad_out_rsc_vld;
  input rec_quad_out_rsc_rdy;
  output [46:0] closest_so_far_out_rsc_dat;
  output closest_so_far_out_rsc_vld;
  input closest_so_far_out_rsc_rdy;


  // Interconnect Declarations
  wire [33:0] mult_run_mul_cmp_a;
  wire [46:0] mult_run_mul_cmp_b;
  wire mult_run_mul_cmp_en;
  wire [74:0] mult_run_mul_cmp_z;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_b;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_1_b;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_2_b;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_3_b;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_4_b;
  wire [24:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_a;
  wire [55:0] quadInters_qnorm_rorig_run_mul_1_cmp_5_b;
  wire [25:0] quadInters_denom_dot_run_mul_2_cmp_a;
  wire [33:0] quadInters_denom_dot_run_mul_2_cmp_b;
  wire [25:0] quadInters_denom_dot_run_mul_2_cmp_1_a;
  wire [33:0] quadInters_denom_dot_run_mul_2_cmp_1_b;
  wire [25:0] quadInters_denom_dot_run_mul_1_cmp_a;
  wire [33:0] quadInters_denom_dot_run_mul_1_cmp_b;


  // Interconnect Declarations for Component Instantiations 
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_b));
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_1_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_1_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_1_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_1_b));
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_2_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_2_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_2_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_2_b));
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_3_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_3_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_3_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_3_b));
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_4_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_4_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_4_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_4_b));
  wire [61:0] nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_5_z;
  assign nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_5_z = conv_u2u_81_62($signed(quadInters_qnorm_rorig_run_mul_1_cmp_5_a)
      * $signed(quadInters_qnorm_rorig_run_mul_1_cmp_5_b));
  wire [57:0] nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_z;
  assign nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_z = conv_u2u_60_58($signed(quadInters_denom_dot_run_mul_2_cmp_a)
      * $signed(quadInters_denom_dot_run_mul_2_cmp_b));
  wire [57:0] nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_1_z;
  assign nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_1_z = conv_u2u_60_58($signed(quadInters_denom_dot_run_mul_2_cmp_1_a)
      * $signed(quadInters_denom_dot_run_mul_2_cmp_1_b));
  wire [59:0] nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_1_cmp_z;
  assign nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_1_cmp_z = conv_u2u_60_60($signed(quadInters_denom_dot_run_mul_1_cmp_a)
      * $signed(quadInters_denom_dot_run_mul_1_cmp_b));
  mgc_mul_pipe #(.width_a(32'sd34),
  .signd_a(32'sd1),
  .width_b(32'sd47),
  .signd_b(32'sd1),
  .width_z(32'sd75),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_run_mul_cmp (
      .a(mult_run_mul_cmp_a),
      .b(mult_run_mul_cmp_b),
      .clk(clk),
      .en(mult_run_mul_cmp_en),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .z(mult_run_mul_cmp_z)
    );
  IntersecLoop_hit IntersecLoop_hit_inst (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsc_dat(quads_rsc_dat),
      .quads_rsc_vld(quads_rsc_vld),
      .quads_rsc_rdy(quads_rsc_rdy),
      .ray_temp_in_rsc_dat(ray_temp_in_rsc_dat),
      .ray_temp_in_rsc_vld(ray_temp_in_rsc_vld),
      .ray_temp_in_rsc_rdy(ray_temp_in_rsc_rdy),
      .quad_max_in_rsc_dat(quad_max_in_rsc_dat),
      .quad_max_in_rsc_vld(quad_max_in_rsc_vld),
      .quad_max_in_rsc_rdy(quad_max_in_rsc_rdy),
      .quad_hit_anything_out_rsc_dat(quad_hit_anything_out_rsc_dat),
      .quad_hit_anything_out_rsc_vld(quad_hit_anything_out_rsc_vld),
      .quad_hit_anything_out_rsc_rdy(quad_hit_anything_out_rsc_rdy),
      .rec_quad_out_rsc_dat(rec_quad_out_rsc_dat),
      .rec_quad_out_rsc_vld(rec_quad_out_rsc_vld),
      .rec_quad_out_rsc_rdy(rec_quad_out_rsc_rdy),
      .closest_so_far_out_rsc_dat(closest_so_far_out_rsc_dat),
      .closest_so_far_out_rsc_vld(closest_so_far_out_rsc_vld),
      .closest_so_far_out_rsc_rdy(closest_so_far_out_rsc_rdy),
      .mult_run_mul_cmp_a(mult_run_mul_cmp_a),
      .mult_run_mul_cmp_b(mult_run_mul_cmp_b),
      .mult_run_mul_cmp_en(mult_run_mul_cmp_en),
      .mult_run_mul_cmp_z(mult_run_mul_cmp_z),
      .quadInters_qnorm_rorig_run_mul_1_cmp_a(quadInters_qnorm_rorig_run_mul_1_cmp_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_b(quadInters_qnorm_rorig_run_mul_1_cmp_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_z[61:0]),
      .quadInters_qnorm_rorig_run_mul_1_cmp_1_a(quadInters_qnorm_rorig_run_mul_1_cmp_1_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_1_b(quadInters_qnorm_rorig_run_mul_1_cmp_1_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_1_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_1_z[61:0]),
      .quadInters_qnorm_rorig_run_mul_1_cmp_2_a(quadInters_qnorm_rorig_run_mul_1_cmp_2_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_2_b(quadInters_qnorm_rorig_run_mul_1_cmp_2_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_2_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_2_z[61:0]),
      .quadInters_qnorm_rorig_run_mul_1_cmp_3_a(quadInters_qnorm_rorig_run_mul_1_cmp_3_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_3_b(quadInters_qnorm_rorig_run_mul_1_cmp_3_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_3_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_3_z[61:0]),
      .quadInters_qnorm_rorig_run_mul_1_cmp_4_a(quadInters_qnorm_rorig_run_mul_1_cmp_4_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_4_b(quadInters_qnorm_rorig_run_mul_1_cmp_4_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_4_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_4_z[61:0]),
      .quadInters_qnorm_rorig_run_mul_1_cmp_5_a(quadInters_qnorm_rorig_run_mul_1_cmp_5_a),
      .quadInters_qnorm_rorig_run_mul_1_cmp_5_b(quadInters_qnorm_rorig_run_mul_1_cmp_5_b),
      .quadInters_qnorm_rorig_run_mul_1_cmp_5_z(nl_IntersecLoop_hit_inst_quadInters_qnorm_rorig_run_mul_1_cmp_5_z[61:0]),
      .quadInters_denom_dot_run_mul_2_cmp_a(quadInters_denom_dot_run_mul_2_cmp_a),
      .quadInters_denom_dot_run_mul_2_cmp_b(quadInters_denom_dot_run_mul_2_cmp_b),
      .quadInters_denom_dot_run_mul_2_cmp_z(nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_z[57:0]),
      .quadInters_denom_dot_run_mul_2_cmp_1_a(quadInters_denom_dot_run_mul_2_cmp_1_a),
      .quadInters_denom_dot_run_mul_2_cmp_1_b(quadInters_denom_dot_run_mul_2_cmp_1_b),
      .quadInters_denom_dot_run_mul_2_cmp_1_z(nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_2_cmp_1_z[57:0]),
      .quadInters_denom_dot_run_mul_1_cmp_a(quadInters_denom_dot_run_mul_1_cmp_a),
      .quadInters_denom_dot_run_mul_1_cmp_b(quadInters_denom_dot_run_mul_1_cmp_b),
      .quadInters_denom_dot_run_mul_1_cmp_z(nl_IntersecLoop_hit_inst_quadInters_denom_dot_run_mul_1_cmp_z[59:0])
    );

  function automatic [57:0] conv_u2u_60_58 ;
    input [59:0]  vector ;
  begin
    conv_u2u_60_58 = vector[57:0];
  end
  endfunction


  function automatic [59:0] conv_u2u_60_60 ;
    input [59:0]  vector ;
  begin
    conv_u2u_60_60 = vector;
  end
  endfunction


  function automatic [61:0] conv_u2u_81_62 ;
    input [80:0]  vector ;
  begin
    conv_u2u_81_62 = vector[61:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    WorldHit
// ------------------------------------------------------------------


module WorldHit (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld,
      attenuation_chan_in_rsc_rdy, accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld,
      accumalated_color_chan_in_rsc_rdy, quad_hit_anything_outone_rsc_dat, quad_hit_anything_outone_rsc_vld,
      quad_hit_anything_outone_rsc_rdy, quad_hit_anything_outtwo_rsc_dat, quad_hit_anything_outtwo_rsc_vld,
      quad_hit_anything_outtwo_rsc_rdy, rec_quad_outone_rsc_dat, rec_quad_outone_rsc_vld,
      rec_quad_outone_rsc_rdy, rec_quad_outtwo_rsc_dat, rec_quad_outtwo_rsc_vld,
      rec_quad_outtwo_rsc_rdy, closest_so_far_outone_rsc_dat, closest_so_far_outone_rsc_vld,
      closest_so_far_outone_rsc_rdy, closest_so_far_outtwo_rsc_dat, closest_so_far_outtwo_rsc_vld,
      closest_so_far_outtwo_rsc_rdy, attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld,
      attenuation_chan_out_rsc_rdy, accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld,
      accumalated_color_out_rsc_rdy, hit_out_rsc_dat, hit_out_rsc_vld, hit_out_rsc_rdy,
      ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, isHit_rsc_dat, isHit_rsc_vld,
      isHit_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input quad_hit_anything_outone_rsc_dat;
  input quad_hit_anything_outone_rsc_vld;
  output quad_hit_anything_outone_rsc_rdy;
  input quad_hit_anything_outtwo_rsc_dat;
  input quad_hit_anything_outtwo_rsc_vld;
  output quad_hit_anything_outtwo_rsc_rdy;
  input [225:0] rec_quad_outone_rsc_dat;
  input rec_quad_outone_rsc_vld;
  output rec_quad_outone_rsc_rdy;
  input [225:0] rec_quad_outtwo_rsc_dat;
  input rec_quad_outtwo_rsc_vld;
  output rec_quad_outtwo_rsc_rdy;
  input [46:0] closest_so_far_outone_rsc_dat;
  input closest_so_far_outone_rsc_vld;
  output closest_so_far_outone_rsc_rdy;
  input [46:0] closest_so_far_outtwo_rsc_dat;
  input closest_so_far_outtwo_rsc_vld;
  output closest_so_far_outtwo_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [225:0] hit_out_rsc_dat;
  output hit_out_rsc_vld;
  input hit_out_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  output isHit_rsc_dat;
  output isHit_rsc_vld;
  input isHit_rsc_rdy;


  // Interconnect Declarations
  wire [26:0] else_mul_cmp_a;
  wire [26:0] else_mul_cmp_b;


  // Interconnect Declarations for Component Instantiations 
  wire [48:0] nl_WorldHit_hit_inst_else_mul_cmp_z;
  assign nl_WorldHit_hit_inst_else_mul_cmp_z = conv_u2u_54_49(else_mul_cmp_a * else_mul_cmp_b);
  WorldHit_hit WorldHit_hit_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .quad_hit_anything_outone_rsc_dat(quad_hit_anything_outone_rsc_dat),
      .quad_hit_anything_outone_rsc_vld(quad_hit_anything_outone_rsc_vld),
      .quad_hit_anything_outone_rsc_rdy(quad_hit_anything_outone_rsc_rdy),
      .quad_hit_anything_outtwo_rsc_dat(quad_hit_anything_outtwo_rsc_dat),
      .quad_hit_anything_outtwo_rsc_vld(quad_hit_anything_outtwo_rsc_vld),
      .quad_hit_anything_outtwo_rsc_rdy(quad_hit_anything_outtwo_rsc_rdy),
      .rec_quad_outone_rsc_dat(rec_quad_outone_rsc_dat),
      .rec_quad_outone_rsc_vld(rec_quad_outone_rsc_vld),
      .rec_quad_outone_rsc_rdy(rec_quad_outone_rsc_rdy),
      .rec_quad_outtwo_rsc_dat(rec_quad_outtwo_rsc_dat),
      .rec_quad_outtwo_rsc_vld(rec_quad_outtwo_rsc_vld),
      .rec_quad_outtwo_rsc_rdy(rec_quad_outtwo_rsc_rdy),
      .closest_so_far_outone_rsc_dat(closest_so_far_outone_rsc_dat),
      .closest_so_far_outone_rsc_vld(closest_so_far_outone_rsc_vld),
      .closest_so_far_outone_rsc_rdy(closest_so_far_outone_rsc_rdy),
      .closest_so_far_outtwo_rsc_dat(closest_so_far_outtwo_rsc_dat),
      .closest_so_far_outtwo_rsc_vld(closest_so_far_outtwo_rsc_vld),
      .closest_so_far_outtwo_rsc_rdy(closest_so_far_outtwo_rsc_rdy),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .hit_out_rsc_dat(hit_out_rsc_dat),
      .hit_out_rsc_vld(hit_out_rsc_vld),
      .hit_out_rsc_rdy(hit_out_rsc_rdy),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .isHit_rsc_dat(isHit_rsc_dat),
      .isHit_rsc_vld(isHit_rsc_vld),
      .isHit_rsc_rdy(isHit_rsc_rdy),
      .else_mul_cmp_a(else_mul_cmp_a),
      .else_mul_cmp_b(else_mul_cmp_b),
      .else_mul_cmp_z(nl_WorldHit_hit_inst_else_mul_cmp_z[48:0])
    );

  function automatic [48:0] conv_u2u_54_49 ;
    input [53:0]  vector ;
  begin
    conv_u2u_54_49 = vector[48:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MaterialScatter
// ------------------------------------------------------------------


module MaterialScatter (
  clk, arst_n, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy, hit_in_rsc_dat, hit_in_rsc_vld,
      hit_in_rsc_rdy, attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld, accumalated_color_chan_in_rsc_rdy,
      isHit_rsc_dat, isHit_rsc_vld, isHit_rsc_rdy, attenuation_chan_out_rsc_dat,
      attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy, accumalated_color_out_rsc_dat,
      accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy, ray_out_rsc_dat,
      ray_out_rsc_vld, ray_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [225:0] hit_in_rsc_dat;
  input hit_in_rsc_vld;
  output hit_in_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  input isHit_rsc_dat;
  input isHit_rsc_vld;
  output isHit_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;


  // Interconnect Declarations
  wire [35:0] lambertianScatter_rand_unit_run_xs_mul_cmp_a;
  wire [35:0] lambertianScatter_rand_unit_run_xs_mul_cmp_b;
  wire lambertianScatter_rand_unit_run_xs_mul_cmp_en;
  wire [65:0] lambertianScatter_rand_unit_run_xs_mul_cmp_z;
  wire [26:0] else_if_mul_cmp_a;
  wire [26:0] else_if_mul_cmp_b;


  // Interconnect Declarations for Component Instantiations 
  wire [48:0] nl_MaterialScatter_scatter_inst_else_if_mul_cmp_z;
  assign nl_MaterialScatter_scatter_inst_else_if_mul_cmp_z = conv_u2u_54_49(else_if_mul_cmp_a
      * else_if_mul_cmp_b);
  mgc_mul_pipe #(.width_a(32'sd36),
  .signd_a(32'sd1),
  .width_b(32'sd36),
  .signd_b(32'sd1),
  .width_z(32'sd66),
  .clock_edge(32'sd1),
  .enable_active(32'sd0),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd0),
  .stages(32'sd2),
  .n_inreg(32'sd0)) lambertianScatter_rand_unit_run_xs_mul_cmp (
      .a(lambertianScatter_rand_unit_run_xs_mul_cmp_a),
      .b(lambertianScatter_rand_unit_run_xs_mul_cmp_b),
      .clk(clk),
      .en(lambertianScatter_rand_unit_run_xs_mul_cmp_en),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .z(lambertianScatter_rand_unit_run_xs_mul_cmp_z)
    );
  MaterialScatter_scatter MaterialScatter_scatter_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy),
      .hit_in_rsc_dat(hit_in_rsc_dat),
      .hit_in_rsc_vld(hit_in_rsc_vld),
      .hit_in_rsc_rdy(hit_in_rsc_rdy),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy),
      .isHit_rsc_dat(isHit_rsc_dat),
      .isHit_rsc_vld(isHit_rsc_vld),
      .isHit_rsc_rdy(isHit_rsc_rdy),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_a(lambertianScatter_rand_unit_run_xs_mul_cmp_a),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_b(lambertianScatter_rand_unit_run_xs_mul_cmp_b),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_en(lambertianScatter_rand_unit_run_xs_mul_cmp_en),
      .lambertianScatter_rand_unit_run_xs_mul_cmp_z(lambertianScatter_rand_unit_run_xs_mul_cmp_z),
      .else_if_mul_cmp_a(else_if_mul_cmp_a),
      .else_if_mul_cmp_b(else_if_mul_cmp_b),
      .else_if_mul_cmp_z(nl_MaterialScatter_scatter_inst_else_if_mul_cmp_z[48:0])
    );

  function automatic [48:0] conv_u2u_54_49 ;
    input [53:0]  vector ;
  begin
    conv_u2u_54_49 = vector[48:0];
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderFeedbackController
// ------------------------------------------------------------------


module ShaderFeedbackController (
  clk, arst_n, ray_chan_in_rsc_dat, ray_chan_in_rsc_vld, ray_chan_in_rsc_rdy, ray_scattered_chan_rsc_dat,
      ray_scattered_chan_rsc_vld, ray_scattered_chan_rsc_rdy, params_in_rsc_dat,
      params_in_rsc_vld, params_in_rsc_rdy, color_chan_in_rsc_dat, color_chan_in_rsc_vld,
      color_chan_in_rsc_rdy, atten_chan_in_rsc_dat, atten_chan_in_rsc_vld, atten_chan_in_rsc_rdy,
      ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy, params_out_rsc_dat, params_out_rsc_vld,
      params_out_rsc_rdy, color_chan_out_rsc_dat, color_chan_out_rsc_vld, color_chan_out_rsc_rdy,
      atten_chan_out_rsc_dat, atten_chan_out_rsc_vld, atten_chan_out_rsc_rdy, output_pxl_serial_rsc_dat,
      output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] ray_chan_in_rsc_dat;
  input ray_chan_in_rsc_vld;
  output ray_chan_in_rsc_rdy;
  input [165:0] ray_scattered_chan_rsc_dat;
  input ray_scattered_chan_rsc_vld;
  output ray_scattered_chan_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [80:0] color_chan_in_rsc_dat;
  input color_chan_in_rsc_vld;
  output color_chan_in_rsc_rdy;
  input [80:0] atten_chan_in_rsc_dat;
  input atten_chan_in_rsc_vld;
  output atten_chan_in_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;
  output [92:0] params_out_rsc_dat;
  output params_out_rsc_vld;
  input params_out_rsc_rdy;
  output [80:0] color_chan_out_rsc_dat;
  output color_chan_out_rsc_vld;
  input color_chan_out_rsc_rdy;
  output [80:0] atten_chan_out_rsc_dat;
  output atten_chan_out_rsc_vld;
  input atten_chan_out_rsc_rdy;
  output [80:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ShaderFeedbackController_run ShaderFeedbackController_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ray_chan_in_rsc_dat(ray_chan_in_rsc_dat),
      .ray_chan_in_rsc_vld(ray_chan_in_rsc_vld),
      .ray_chan_in_rsc_rdy(ray_chan_in_rsc_rdy),
      .ray_scattered_chan_rsc_dat(ray_scattered_chan_rsc_dat),
      .ray_scattered_chan_rsc_vld(ray_scattered_chan_rsc_vld),
      .ray_scattered_chan_rsc_rdy(ray_scattered_chan_rsc_rdy),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy),
      .color_chan_in_rsc_dat(color_chan_in_rsc_dat),
      .color_chan_in_rsc_vld(color_chan_in_rsc_vld),
      .color_chan_in_rsc_rdy(color_chan_in_rsc_rdy),
      .atten_chan_in_rsc_dat(atten_chan_in_rsc_dat),
      .atten_chan_in_rsc_vld(atten_chan_in_rsc_vld),
      .atten_chan_in_rsc_rdy(atten_chan_in_rsc_rdy),
      .ray_out_rsc_dat(ray_out_rsc_dat),
      .ray_out_rsc_vld(ray_out_rsc_vld),
      .ray_out_rsc_rdy(ray_out_rsc_rdy),
      .params_out_rsc_dat(params_out_rsc_dat),
      .params_out_rsc_vld(params_out_rsc_vld),
      .params_out_rsc_rdy(params_out_rsc_rdy),
      .color_chan_out_rsc_dat(color_chan_out_rsc_dat),
      .color_chan_out_rsc_vld(color_chan_out_rsc_vld),
      .color_chan_out_rsc_rdy(color_chan_out_rsc_rdy),
      .atten_chan_out_rsc_dat(atten_chan_out_rsc_dat),
      .atten_chan_out_rsc_vld(atten_chan_out_rsc_vld),
      .atten_chan_out_rsc_rdy(atten_chan_out_rsc_rdy),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    RayCollector
// ------------------------------------------------------------------


module RayCollector (
  clk, arst_n, rayIn_rsc_dat, rayIn_rsc_vld, rayIn_rsc_rdy, paramsIn_rsc_dat, paramsIn_rsc_vld,
      paramsIn_rsc_rdy, paramsOut_rsc_dat, paramsOut_rsc_vld, paramsOut_rsc_rdy,
      rayOut_rsc_dat, rayOut_rsc_vld, rayOut_rsc_rdy
);
  input clk;
  input arst_n;
  input [165:0] rayIn_rsc_dat;
  input rayIn_rsc_vld;
  output rayIn_rsc_rdy;
  input [92:0] paramsIn_rsc_dat;
  input paramsIn_rsc_vld;
  output paramsIn_rsc_rdy;
  output [92:0] paramsOut_rsc_dat;
  output paramsOut_rsc_vld;
  input paramsOut_rsc_rdy;
  output [165:0] rayOut_rsc_dat;
  output rayOut_rsc_vld;
  input rayOut_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  RayCollector_run RayCollector_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .rayIn_rsc_dat(rayIn_rsc_dat),
      .rayIn_rsc_vld(rayIn_rsc_vld),
      .rayIn_rsc_rdy(rayIn_rsc_rdy),
      .paramsIn_rsc_dat(paramsIn_rsc_dat),
      .paramsIn_rsc_vld(paramsIn_rsc_vld),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy),
      .paramsOut_rsc_dat(paramsOut_rsc_dat),
      .paramsOut_rsc_vld(paramsOut_rsc_vld),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy),
      .rayOut_rsc_dat(rayOut_rsc_dat),
      .rayOut_rsc_vld(rayOut_rsc_vld),
      .rayOut_rsc_rdy(rayOut_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    PixelAccumulator
// ------------------------------------------------------------------


module PixelAccumulator (
  clk, arst_n, accumulator_parms_rsc_dat, accumulator_parms_rsc_vld, accumulator_parms_rsc_rdy,
      pxl_sample_rsc_dat, pxl_sample_rsc_vld, pxl_sample_rsc_rdy, output_pxl_serial_rsc_dat,
      output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [419:0] accumulator_parms_rsc_dat;
  input accumulator_parms_rsc_vld;
  output accumulator_parms_rsc_rdy;
  input [80:0] pxl_sample_rsc_dat;
  input pxl_sample_rsc_vld;
  output pxl_sample_rsc_rdy;
  output [23:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  PixelAccumulator_run PixelAccumulator_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .accumulator_parms_rsc_dat(accumulator_parms_rsc_dat),
      .accumulator_parms_rsc_vld(accumulator_parms_rsc_vld),
      .accumulator_parms_rsc_rdy(accumulator_parms_rsc_rdy),
      .pxl_sample_rsc_dat(pxl_sample_rsc_dat),
      .pxl_sample_rsc_vld(pxl_sample_rsc_vld),
      .pxl_sample_rsc_rdy(pxl_sample_rsc_rdy),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Shader
// ------------------------------------------------------------------


module Shader (
  clk, arst_n, params_in_rsc_dat, params_in_rsc_vld, params_in_rsc_rdy, quad_in_rsc_dat,
      quad_in_rsc_vld, quad_in_rsc_rdy, ray_in_rsc_dat, ray_in_rsc_vld, ray_in_rsc_rdy,
      attenuation_chan_in_rsc_dat, attenuation_chan_in_rsc_vld, attenuation_chan_in_rsc_rdy,
      accumalated_color_chan_in_rsc_dat, accumalated_color_chan_in_rsc_vld, accumalated_color_chan_in_rsc_rdy,
      attenuation_chan_out_rsc_dat, attenuation_chan_out_rsc_vld, attenuation_chan_out_rsc_rdy,
      accumalated_color_out_rsc_dat, accumalated_color_out_rsc_vld, accumalated_color_out_rsc_rdy,
      ray_out_rsc_dat, ray_out_rsc_vld, ray_out_rsc_rdy
);
  input clk;
  input arst_n;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  input [376:0] quad_in_rsc_dat;
  input quad_in_rsc_vld;
  output quad_in_rsc_rdy;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [80:0] attenuation_chan_in_rsc_dat;
  input attenuation_chan_in_rsc_vld;
  output attenuation_chan_in_rsc_rdy;
  input [80:0] accumalated_color_chan_in_rsc_dat;
  input accumalated_color_chan_in_rsc_vld;
  output accumalated_color_chan_in_rsc_rdy;
  output [80:0] attenuation_chan_out_rsc_dat;
  output attenuation_chan_out_rsc_vld;
  input attenuation_chan_out_rsc_rdy;
  output [80:0] accumalated_color_out_rsc_dat;
  output accumalated_color_out_rsc_vld;
  input accumalated_color_out_rsc_rdy;
  output [165:0] ray_out_rsc_dat;
  output ray_out_rsc_vld;
  input ray_out_rsc_rdy;


  // Interconnect Declarations
  wire [80:0] attenuation_chan_out_rsc_dat_nloop_distrib;
  wire attenuation_chan_out_rsc_rdy_nloop_distrib;
  wire [80:0] accumalated_color_out_rsc_dat_nloop_distrib;
  wire accumalated_color_out_rsc_rdy_nloop_distrib;
  wire [165:0] ray_out_loopone_rsc_dat_nloop_distrib;
  wire ray_out_loopone_rsc_rdy_nloop_distrib;
  wire [165:0] ray_out_looptwo_rsc_dat_nloop_distrib;
  wire ray_out_looptwo_rsc_rdy_nloop_distrib;
  wire [165:0] ray_out_worldhit_rsc_dat_nloop_distrib;
  wire ray_out_worldhit_rsc_rdy_nloop_distrib;
  wire [376:0] quad_out_loopone_rsc_dat_nloop_distrib;
  wire quad_out_loopone_rsc_rdy_nloop_distrib;
  wire [376:0] quad_out_looptwo_rsc_dat_nloop_distrib;
  wire quad_out_looptwo_rsc_rdy_nloop_distrib;
  wire [10:0] quad_max_outone_rsc_dat_nloop_distrib;
  wire quad_max_outone_rsc_rdy_nloop_distrib;
  wire [10:0] quad_max_outtwo_rsc_dat_nloop_distrib;
  wire quad_max_outtwo_rsc_rdy_nloop_distrib;
  wire [92:0] params_out_rsc_dat_nloop_distrib;
  wire params_out_rsc_rdy_nloop_distrib;
  wire [376:0] quads_rsc_dat_nintersec_loop_one;
  wire quads_rsc_vld_nintersec_loop_one;
  wire [165:0] ray_temp_in_rsc_dat_nintersec_loop_one;
  wire ray_temp_in_rsc_vld_nintersec_loop_one;
  wire [10:0] quad_max_in_rsc_dat_nintersec_loop_one;
  wire quad_max_in_rsc_vld_nintersec_loop_one;
  wire quad_hit_anything_out_rsc_dat_nintersec_loop_one;
  wire quad_hit_anything_out_rsc_rdy_nintersec_loop_one;
  wire [225:0] rec_quad_out_rsc_dat_nintersec_loop_one;
  wire rec_quad_out_rsc_rdy_nintersec_loop_one;
  wire [46:0] closest_so_far_out_rsc_dat_nintersec_loop_one;
  wire closest_so_far_out_rsc_rdy_nintersec_loop_one;
  wire [376:0] quads_rsc_dat_nintersec_loop_two;
  wire quads_rsc_vld_nintersec_loop_two;
  wire [165:0] ray_temp_in_rsc_dat_nintersec_loop_two;
  wire ray_temp_in_rsc_vld_nintersec_loop_two;
  wire [10:0] quad_max_in_rsc_dat_nintersec_loop_two;
  wire quad_max_in_rsc_vld_nintersec_loop_two;
  wire quad_hit_anything_out_rsc_dat_nintersec_loop_two;
  wire quad_hit_anything_out_rsc_rdy_nintersec_loop_two;
  wire [225:0] rec_quad_out_rsc_dat_nintersec_loop_two;
  wire rec_quad_out_rsc_rdy_nintersec_loop_two;
  wire [46:0] closest_so_far_out_rsc_dat_nintersec_loop_two;
  wire closest_so_far_out_rsc_rdy_nintersec_loop_two;
  wire [165:0] ray_in_rsc_dat_nworldHit;
  wire ray_in_rsc_vld_nworldHit;
  wire [92:0] params_in_rsc_dat_nworldHit;
  wire params_in_rsc_vld_nworldHit;
  wire [80:0] attenuation_chan_in_rsc_dat_nworldHit;
  wire attenuation_chan_in_rsc_vld_nworldHit;
  wire [80:0] accumalated_color_chan_in_rsc_dat_nworldHit;
  wire accumalated_color_chan_in_rsc_vld_nworldHit;
  wire quad_hit_anything_outone_rsc_dat_nworldHit;
  wire quad_hit_anything_outone_rsc_vld_nworldHit;
  wire quad_hit_anything_outtwo_rsc_dat_nworldHit;
  wire quad_hit_anything_outtwo_rsc_vld_nworldHit;
  wire [225:0] rec_quad_outone_rsc_dat_nworldHit;
  wire rec_quad_outone_rsc_vld_nworldHit;
  wire [225:0] rec_quad_outtwo_rsc_dat_nworldHit;
  wire rec_quad_outtwo_rsc_vld_nworldHit;
  wire [46:0] closest_so_far_outone_rsc_dat_nworldHit;
  wire closest_so_far_outone_rsc_vld_nworldHit;
  wire [46:0] closest_so_far_outtwo_rsc_dat_nworldHit;
  wire closest_so_far_outtwo_rsc_vld_nworldHit;
  wire [80:0] attenuation_chan_out_rsc_dat_nworldHit;
  wire attenuation_chan_out_rsc_rdy_nworldHit;
  wire [80:0] accumalated_color_out_rsc_dat_nworldHit;
  wire accumalated_color_out_rsc_rdy_nworldHit;
  wire [225:0] hit_out_rsc_dat_nworldHit;
  wire hit_out_rsc_rdy_nworldHit;
  wire [165:0] ray_out_rsc_dat_nworldHit;
  wire ray_out_rsc_rdy_nworldHit;
  wire isHit_rsc_dat_nworldHit;
  wire isHit_rsc_rdy_nworldHit;
  wire [165:0] ray_in_rsc_dat_nmaterialScatter;
  wire ray_in_rsc_vld_nmaterialScatter;
  wire [225:0] hit_in_rsc_dat_nmaterialScatter;
  wire hit_in_rsc_vld_nmaterialScatter;
  wire [80:0] attenuation_chan_in_rsc_dat_nmaterialScatter;
  wire attenuation_chan_in_rsc_vld_nmaterialScatter;
  wire [80:0] accumalated_color_chan_in_rsc_dat_nmaterialScatter;
  wire accumalated_color_chan_in_rsc_vld_nmaterialScatter;
  wire isHit_rsc_dat_nmaterialScatter;
  wire isHit_rsc_vld_nmaterialScatter;
  wire [80:0] attenuation_chan_out_rsc_dat_nmaterialScatter;
  wire [80:0] accumalated_color_out_rsc_dat_nmaterialScatter;
  wire [165:0] ray_out_rsc_dat_nmaterialScatter;
  wire ray_in_rsc_rdy_nloop_distrib_bud;
  wire params_in_rsc_rdy_nloop_distrib_bud;
  wire quads_rsc_rdy_nloop_distrib_bud;
  wire attenuation_chan_in_rsc_rdy_nloop_distrib_bud;
  wire accumalated_color_chan_in_rsc_rdy_nloop_distrib_bud;
  wire attenuation_chan_out_rsc_vld_nloop_distrib_bud;
  wire attenuation_chan_in_rsc_rdy_nworldHit_bud;
  wire accumalated_color_out_rsc_vld_nloop_distrib_bud;
  wire accumalated_color_chan_in_rsc_rdy_nworldHit_bud;
  wire ray_out_loopone_rsc_vld_nloop_distrib_bud;
  wire ray_temp_in_rsc_rdy_nintersec_loop_one_bud;
  wire ray_out_looptwo_rsc_vld_nloop_distrib_bud;
  wire ray_temp_in_rsc_rdy_nintersec_loop_two_bud;
  wire ray_out_worldhit_rsc_vld_nloop_distrib_bud;
  wire ray_in_rsc_rdy_nworldHit_bud;
  wire quad_out_loopone_rsc_vld_nloop_distrib_bud;
  wire quads_rsc_rdy_nintersec_loop_one_bud;
  wire quad_out_looptwo_rsc_vld_nloop_distrib_bud;
  wire quads_rsc_rdy_nintersec_loop_two_bud;
  wire quad_max_outone_rsc_vld_nloop_distrib_bud;
  wire quad_max_in_rsc_rdy_nintersec_loop_one_bud;
  wire quad_max_outtwo_rsc_vld_nloop_distrib_bud;
  wire quad_max_in_rsc_rdy_nintersec_loop_two_bud;
  wire params_out_rsc_vld_nloop_distrib_bud;
  wire params_in_rsc_rdy_nworldHit_bud;
  wire quad_hit_anything_out_rsc_vld_nintersec_loop_one_bud;
  wire quad_hit_anything_outone_rsc_rdy_nworldHit_bud;
  wire rec_quad_out_rsc_vld_nintersec_loop_one_bud;
  wire rec_quad_outone_rsc_rdy_nworldHit_bud;
  wire closest_so_far_out_rsc_vld_nintersec_loop_one_bud;
  wire closest_so_far_outone_rsc_rdy_nworldHit_bud;
  wire quad_hit_anything_out_rsc_vld_nintersec_loop_two_bud;
  wire quad_hit_anything_outtwo_rsc_rdy_nworldHit_bud;
  wire rec_quad_out_rsc_vld_nintersec_loop_two_bud;
  wire rec_quad_outtwo_rsc_rdy_nworldHit_bud;
  wire closest_so_far_out_rsc_vld_nintersec_loop_two_bud;
  wire closest_so_far_outtwo_rsc_rdy_nworldHit_bud;
  wire attenuation_chan_out_rsc_vld_nworldHit_bud;
  wire attenuation_chan_in_rsc_rdy_nmaterialScatter_bud;
  wire accumalated_color_out_rsc_vld_nworldHit_bud;
  wire accumalated_color_chan_in_rsc_rdy_nmaterialScatter_bud;
  wire hit_out_rsc_vld_nworldHit_bud;
  wire hit_in_rsc_rdy_nmaterialScatter_bud;
  wire ray_out_rsc_vld_nworldHit_bud;
  wire ray_in_rsc_rdy_nmaterialScatter_bud;
  wire isHit_rsc_vld_nworldHit_bud;
  wire isHit_rsc_rdy_nmaterialScatter_bud;
  wire attenuation_chan_out_rsc_vld_nmaterialScatter_bud;
  wire accumalated_color_out_rsc_vld_nmaterialScatter_bud;
  wire ray_out_rsc_vld_nmaterialScatter_bud;
  wire attenuation_chan_to_WorldHit_unc_2;
  wire attenuation_chan_to_WorldHit_idle;
  wire accumalated_color_to_WorldHit_unc_2;
  wire accumalated_color_to_WorldHit_idle;
  wire rayToLoopOne_unc_2;
  wire rayToLoopOne_idle;
  wire rayToLoopTwo_unc_2;
  wire rayToLoopTwo_idle;
  wire rayToWorldHit_unc_2;
  wire rayToWorldHit_idle;
  wire quad_to_loopone_unc_2;
  wire quad_to_loopone_idle;
  wire quad_to_looptwo_unc_2;
  wire quad_to_looptwo_idle;
  wire quad_max_outone_unc_2;
  wire quad_max_outone_idle;
  wire quad_max_outtwo_unc_2;
  wire quad_max_outtwo_idle;
  wire params_to_WorldHit_unc_2;
  wire params_to_WorldHit_idle;
  wire quad_hit_anything_outone_unc_2;
  wire quad_hit_anything_outone_idle;
  wire rec_quad_outone_unc_2;
  wire rec_quad_outone_idle;
  wire closest_so_far_outone_unc_2;
  wire closest_so_far_outone_idle;
  wire quad_hit_anything_outtwo_unc_2;
  wire quad_hit_anything_outtwo_idle;
  wire rec_quad_outtwo_unc_2;
  wire rec_quad_outtwo_idle;
  wire closest_so_far_outtwo_unc_2;
  wire closest_so_far_outtwo_idle;
  wire attenuation_chan_through_unc_2;
  wire attenuation_chan_through_idle;
  wire accumalated_color_through_unc_2;
  wire accumalated_color_through_idle;
  wire worldRec_unc_2;
  wire worldRec_idle;
  wire rayToScatter_unc_2;
  wire rayToScatter_idle;
  wire isWorldHit_unc_2;
  wire isWorldHit_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd97),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) attenuation_chan_to_WorldHit_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(attenuation_chan_out_rsc_rdy_nloop_distrib),
      .din_vld(attenuation_chan_out_rsc_vld_nloop_distrib_bud),
      .din(attenuation_chan_out_rsc_dat_nloop_distrib),
      .dout_rdy(attenuation_chan_in_rsc_rdy_nworldHit_bud),
      .dout_vld(attenuation_chan_in_rsc_vld_nworldHit),
      .dout(attenuation_chan_in_rsc_dat_nworldHit),
      .sz(attenuation_chan_to_WorldHit_unc_2),
      .sz_req(1'b0),
      .is_idle(attenuation_chan_to_WorldHit_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd98),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) accumalated_color_to_WorldHit_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(accumalated_color_out_rsc_rdy_nloop_distrib),
      .din_vld(accumalated_color_out_rsc_vld_nloop_distrib_bud),
      .din(accumalated_color_out_rsc_dat_nloop_distrib),
      .dout_rdy(accumalated_color_chan_in_rsc_rdy_nworldHit_bud),
      .dout_vld(accumalated_color_chan_in_rsc_vld_nworldHit),
      .dout(accumalated_color_chan_in_rsc_dat_nworldHit),
      .sz(accumalated_color_to_WorldHit_unc_2),
      .sz_req(1'b0),
      .is_idle(accumalated_color_to_WorldHit_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd95),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayToLoopOne_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_loopone_rsc_rdy_nloop_distrib),
      .din_vld(ray_out_loopone_rsc_vld_nloop_distrib_bud),
      .din(ray_out_loopone_rsc_dat_nloop_distrib),
      .dout_rdy(ray_temp_in_rsc_rdy_nintersec_loop_one_bud),
      .dout_vld(ray_temp_in_rsc_vld_nintersec_loop_one),
      .dout(ray_temp_in_rsc_dat_nintersec_loop_one),
      .sz(rayToLoopOne_unc_2),
      .sz_req(1'b0),
      .is_idle(rayToLoopOne_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd96),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayToLoopTwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_looptwo_rsc_rdy_nloop_distrib),
      .din_vld(ray_out_looptwo_rsc_vld_nloop_distrib_bud),
      .din(ray_out_looptwo_rsc_dat_nloop_distrib),
      .dout_rdy(ray_temp_in_rsc_rdy_nintersec_loop_two_bud),
      .dout_vld(ray_temp_in_rsc_vld_nintersec_loop_two),
      .dout(ray_temp_in_rsc_dat_nintersec_loop_two),
      .sz(rayToLoopTwo_unc_2),
      .sz_req(1'b0),
      .is_idle(rayToLoopTwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd94),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayToWorldHit_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_worldhit_rsc_rdy_nloop_distrib),
      .din_vld(ray_out_worldhit_rsc_vld_nloop_distrib_bud),
      .din(ray_out_worldhit_rsc_dat_nloop_distrib),
      .dout_rdy(ray_in_rsc_rdy_nworldHit_bud),
      .dout_vld(ray_in_rsc_vld_nworldHit),
      .dout(ray_in_rsc_dat_nworldHit),
      .sz(rayToWorldHit_unc_2),
      .sz_req(1'b0),
      .is_idle(rayToWorldHit_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd99),
  .width(32'sd377),
  .sz_width(32'sd1),
  .fifo_sz(32'sd19),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_to_loopone_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_out_loopone_rsc_rdy_nloop_distrib),
      .din_vld(quad_out_loopone_rsc_vld_nloop_distrib_bud),
      .din(quad_out_loopone_rsc_dat_nloop_distrib),
      .dout_rdy(quads_rsc_rdy_nintersec_loop_one_bud),
      .dout_vld(quads_rsc_vld_nintersec_loop_one),
      .dout(quads_rsc_dat_nintersec_loop_one),
      .sz(quad_to_loopone_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_to_loopone_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd100),
  .width(32'sd377),
  .sz_width(32'sd1),
  .fifo_sz(32'sd19),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_to_looptwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_out_looptwo_rsc_rdy_nloop_distrib),
      .din_vld(quad_out_looptwo_rsc_vld_nloop_distrib_bud),
      .din(quad_out_looptwo_rsc_dat_nloop_distrib),
      .dout_rdy(quads_rsc_rdy_nintersec_loop_two_bud),
      .dout_vld(quads_rsc_vld_nintersec_loop_two),
      .dout(quads_rsc_dat_nintersec_loop_two),
      .sz(quad_to_looptwo_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_to_looptwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd101),
  .width(32'sd11),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_max_outone_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_max_outone_rsc_rdy_nloop_distrib),
      .din_vld(quad_max_outone_rsc_vld_nloop_distrib_bud),
      .din(quad_max_outone_rsc_dat_nloop_distrib),
      .dout_rdy(quad_max_in_rsc_rdy_nintersec_loop_one_bud),
      .dout_vld(quad_max_in_rsc_vld_nintersec_loop_one),
      .dout(quad_max_in_rsc_dat_nintersec_loop_one),
      .sz(quad_max_outone_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_max_outone_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd102),
  .width(32'sd11),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_max_outtwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_max_outtwo_rsc_rdy_nloop_distrib),
      .din_vld(quad_max_outtwo_rsc_vld_nloop_distrib_bud),
      .din(quad_max_outtwo_rsc_dat_nloop_distrib),
      .dout_rdy(quad_max_in_rsc_rdy_nintersec_loop_two_bud),
      .dout_vld(quad_max_in_rsc_vld_nintersec_loop_two),
      .dout(quad_max_in_rsc_dat_nintersec_loop_two),
      .sz(quad_max_outtwo_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_max_outtwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd109),
  .width(32'sd93),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) params_to_WorldHit_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(params_out_rsc_rdy_nloop_distrib),
      .din_vld(params_out_rsc_vld_nloop_distrib_bud),
      .din(params_out_rsc_dat_nloop_distrib),
      .dout_rdy(params_in_rsc_rdy_nworldHit_bud),
      .dout_vld(params_in_rsc_vld_nworldHit),
      .dout(params_in_rsc_dat_nworldHit),
      .sz(params_to_WorldHit_unc_2),
      .sz_req(1'b0),
      .is_idle(params_to_WorldHit_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd103),
  .width(32'sd1),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_hit_anything_outone_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_hit_anything_out_rsc_rdy_nintersec_loop_one),
      .din_vld(quad_hit_anything_out_rsc_vld_nintersec_loop_one_bud),
      .din(quad_hit_anything_out_rsc_dat_nintersec_loop_one),
      .dout_rdy(quad_hit_anything_outone_rsc_rdy_nworldHit_bud),
      .dout_vld(quad_hit_anything_outone_rsc_vld_nworldHit),
      .dout(quad_hit_anything_outone_rsc_dat_nworldHit),
      .sz(quad_hit_anything_outone_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_hit_anything_outone_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd105),
  .width(32'sd226),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rec_quad_outone_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(rec_quad_out_rsc_rdy_nintersec_loop_one),
      .din_vld(rec_quad_out_rsc_vld_nintersec_loop_one_bud),
      .din(rec_quad_out_rsc_dat_nintersec_loop_one),
      .dout_rdy(rec_quad_outone_rsc_rdy_nworldHit_bud),
      .dout_vld(rec_quad_outone_rsc_vld_nworldHit),
      .dout(rec_quad_outone_rsc_dat_nworldHit),
      .sz(rec_quad_outone_unc_2),
      .sz_req(1'b0),
      .is_idle(rec_quad_outone_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd107),
  .width(32'sd47),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) closest_so_far_outone_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(closest_so_far_out_rsc_rdy_nintersec_loop_one),
      .din_vld(closest_so_far_out_rsc_vld_nintersec_loop_one_bud),
      .din(closest_so_far_out_rsc_dat_nintersec_loop_one),
      .dout_rdy(closest_so_far_outone_rsc_rdy_nworldHit_bud),
      .dout_vld(closest_so_far_outone_rsc_vld_nworldHit),
      .dout(closest_so_far_outone_rsc_dat_nworldHit),
      .sz(closest_so_far_outone_unc_2),
      .sz_req(1'b0),
      .is_idle(closest_so_far_outone_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd104),
  .width(32'sd1),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_hit_anything_outtwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_hit_anything_out_rsc_rdy_nintersec_loop_two),
      .din_vld(quad_hit_anything_out_rsc_vld_nintersec_loop_two_bud),
      .din(quad_hit_anything_out_rsc_dat_nintersec_loop_two),
      .dout_rdy(quad_hit_anything_outtwo_rsc_rdy_nworldHit_bud),
      .dout_vld(quad_hit_anything_outtwo_rsc_vld_nworldHit),
      .dout(quad_hit_anything_outtwo_rsc_dat_nworldHit),
      .sz(quad_hit_anything_outtwo_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_hit_anything_outtwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd106),
  .width(32'sd226),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rec_quad_outtwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(rec_quad_out_rsc_rdy_nintersec_loop_two),
      .din_vld(rec_quad_out_rsc_vld_nintersec_loop_two_bud),
      .din(rec_quad_out_rsc_dat_nintersec_loop_two),
      .dout_rdy(rec_quad_outtwo_rsc_rdy_nworldHit_bud),
      .dout_vld(rec_quad_outtwo_rsc_vld_nworldHit),
      .dout(rec_quad_outtwo_rsc_dat_nworldHit),
      .sz(rec_quad_outtwo_unc_2),
      .sz_req(1'b0),
      .is_idle(rec_quad_outtwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd108),
  .width(32'sd47),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) closest_so_far_outtwo_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(closest_so_far_out_rsc_rdy_nintersec_loop_two),
      .din_vld(closest_so_far_out_rsc_vld_nintersec_loop_two_bud),
      .din(closest_so_far_out_rsc_dat_nintersec_loop_two),
      .dout_rdy(closest_so_far_outtwo_rsc_rdy_nworldHit_bud),
      .dout_vld(closest_so_far_outtwo_rsc_vld_nworldHit),
      .dout(closest_so_far_outtwo_rsc_dat_nworldHit),
      .sz(closest_so_far_outtwo_unc_2),
      .sz_req(1'b0),
      .is_idle(closest_so_far_outtwo_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd111),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) attenuation_chan_through_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(attenuation_chan_out_rsc_rdy_nworldHit),
      .din_vld(attenuation_chan_out_rsc_vld_nworldHit_bud),
      .din(attenuation_chan_out_rsc_dat_nworldHit),
      .dout_rdy(attenuation_chan_in_rsc_rdy_nmaterialScatter_bud),
      .dout_vld(attenuation_chan_in_rsc_vld_nmaterialScatter),
      .dout(attenuation_chan_in_rsc_dat_nmaterialScatter),
      .sz(attenuation_chan_through_unc_2),
      .sz_req(1'b0),
      .is_idle(attenuation_chan_through_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd112),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) accumalated_color_through_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(accumalated_color_out_rsc_rdy_nworldHit),
      .din_vld(accumalated_color_out_rsc_vld_nworldHit_bud),
      .din(accumalated_color_out_rsc_dat_nworldHit),
      .dout_rdy(accumalated_color_chan_in_rsc_rdy_nmaterialScatter_bud),
      .dout_vld(accumalated_color_chan_in_rsc_vld_nmaterialScatter),
      .dout(accumalated_color_chan_in_rsc_dat_nmaterialScatter),
      .sz(accumalated_color_through_unc_2),
      .sz_req(1'b0),
      .is_idle(accumalated_color_through_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd114),
  .width(32'sd226),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) worldRec_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(hit_out_rsc_rdy_nworldHit),
      .din_vld(hit_out_rsc_vld_nworldHit_bud),
      .din(hit_out_rsc_dat_nworldHit),
      .dout_rdy(hit_in_rsc_rdy_nmaterialScatter_bud),
      .dout_vld(hit_in_rsc_vld_nmaterialScatter),
      .dout(hit_in_rsc_dat_nmaterialScatter),
      .sz(worldRec_unc_2),
      .sz_req(1'b0),
      .is_idle(worldRec_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd110),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayToScatter_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_rsc_rdy_nworldHit),
      .din_vld(ray_out_rsc_vld_nworldHit_bud),
      .din(ray_out_rsc_dat_nworldHit),
      .dout_rdy(ray_in_rsc_rdy_nmaterialScatter_bud),
      .dout_vld(ray_in_rsc_vld_nmaterialScatter),
      .dout(ray_in_rsc_dat_nmaterialScatter),
      .sz(rayToScatter_unc_2),
      .sz_req(1'b0),
      .is_idle(rayToScatter_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd113),
  .width(32'sd1),
  .sz_width(32'sd1),
  .fifo_sz(32'sd3),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) isWorldHit_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(isHit_rsc_rdy_nworldHit),
      .din_vld(isHit_rsc_vld_nworldHit_bud),
      .din(isHit_rsc_dat_nworldHit),
      .dout_rdy(isHit_rsc_rdy_nmaterialScatter_bud),
      .dout_vld(isHit_rsc_vld_nmaterialScatter),
      .dout(isHit_rsc_dat_nmaterialScatter),
      .sz(isWorldHit_unc_2),
      .sz_req(1'b0),
      .is_idle(isWorldHit_idle)
    );
  LoopDistrib loop_distrib (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat),
      .ray_in_rsc_vld(ray_in_rsc_vld),
      .ray_in_rsc_rdy(ray_in_rsc_rdy_nloop_distrib_bud),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy_nloop_distrib_bud),
      .quads_rsc_dat(quad_in_rsc_dat),
      .quads_rsc_vld(quad_in_rsc_vld),
      .quads_rsc_rdy(quads_rsc_rdy_nloop_distrib_bud),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy_nloop_distrib_bud),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy_nloop_distrib_bud),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat_nloop_distrib),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld_nloop_distrib_bud),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy_nloop_distrib),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat_nloop_distrib),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld_nloop_distrib_bud),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy_nloop_distrib),
      .ray_out_loopone_rsc_dat(ray_out_loopone_rsc_dat_nloop_distrib),
      .ray_out_loopone_rsc_vld(ray_out_loopone_rsc_vld_nloop_distrib_bud),
      .ray_out_loopone_rsc_rdy(ray_out_loopone_rsc_rdy_nloop_distrib),
      .ray_out_looptwo_rsc_dat(ray_out_looptwo_rsc_dat_nloop_distrib),
      .ray_out_looptwo_rsc_vld(ray_out_looptwo_rsc_vld_nloop_distrib_bud),
      .ray_out_looptwo_rsc_rdy(ray_out_looptwo_rsc_rdy_nloop_distrib),
      .ray_out_worldhit_rsc_dat(ray_out_worldhit_rsc_dat_nloop_distrib),
      .ray_out_worldhit_rsc_vld(ray_out_worldhit_rsc_vld_nloop_distrib_bud),
      .ray_out_worldhit_rsc_rdy(ray_out_worldhit_rsc_rdy_nloop_distrib),
      .quad_out_loopone_rsc_dat(quad_out_loopone_rsc_dat_nloop_distrib),
      .quad_out_loopone_rsc_vld(quad_out_loopone_rsc_vld_nloop_distrib_bud),
      .quad_out_loopone_rsc_rdy(quad_out_loopone_rsc_rdy_nloop_distrib),
      .quad_out_looptwo_rsc_dat(quad_out_looptwo_rsc_dat_nloop_distrib),
      .quad_out_looptwo_rsc_vld(quad_out_looptwo_rsc_vld_nloop_distrib_bud),
      .quad_out_looptwo_rsc_rdy(quad_out_looptwo_rsc_rdy_nloop_distrib),
      .quad_max_outone_rsc_dat(quad_max_outone_rsc_dat_nloop_distrib),
      .quad_max_outone_rsc_vld(quad_max_outone_rsc_vld_nloop_distrib_bud),
      .quad_max_outone_rsc_rdy(quad_max_outone_rsc_rdy_nloop_distrib),
      .quad_max_outtwo_rsc_dat(quad_max_outtwo_rsc_dat_nloop_distrib),
      .quad_max_outtwo_rsc_vld(quad_max_outtwo_rsc_vld_nloop_distrib_bud),
      .quad_max_outtwo_rsc_rdy(quad_max_outtwo_rsc_rdy_nloop_distrib),
      .params_out_rsc_dat(params_out_rsc_dat_nloop_distrib),
      .params_out_rsc_vld(params_out_rsc_vld_nloop_distrib_bud),
      .params_out_rsc_rdy(params_out_rsc_rdy_nloop_distrib)
    );
  IntersecLoop intersec_loop_one (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsc_dat(quads_rsc_dat_nintersec_loop_one),
      .quads_rsc_vld(quads_rsc_vld_nintersec_loop_one),
      .quads_rsc_rdy(quads_rsc_rdy_nintersec_loop_one_bud),
      .ray_temp_in_rsc_dat(ray_temp_in_rsc_dat_nintersec_loop_one),
      .ray_temp_in_rsc_vld(ray_temp_in_rsc_vld_nintersec_loop_one),
      .ray_temp_in_rsc_rdy(ray_temp_in_rsc_rdy_nintersec_loop_one_bud),
      .quad_max_in_rsc_dat(quad_max_in_rsc_dat_nintersec_loop_one),
      .quad_max_in_rsc_vld(quad_max_in_rsc_vld_nintersec_loop_one),
      .quad_max_in_rsc_rdy(quad_max_in_rsc_rdy_nintersec_loop_one_bud),
      .quad_hit_anything_out_rsc_dat(quad_hit_anything_out_rsc_dat_nintersec_loop_one),
      .quad_hit_anything_out_rsc_vld(quad_hit_anything_out_rsc_vld_nintersec_loop_one_bud),
      .quad_hit_anything_out_rsc_rdy(quad_hit_anything_out_rsc_rdy_nintersec_loop_one),
      .rec_quad_out_rsc_dat(rec_quad_out_rsc_dat_nintersec_loop_one),
      .rec_quad_out_rsc_vld(rec_quad_out_rsc_vld_nintersec_loop_one_bud),
      .rec_quad_out_rsc_rdy(rec_quad_out_rsc_rdy_nintersec_loop_one),
      .closest_so_far_out_rsc_dat(closest_so_far_out_rsc_dat_nintersec_loop_one),
      .closest_so_far_out_rsc_vld(closest_so_far_out_rsc_vld_nintersec_loop_one_bud),
      .closest_so_far_out_rsc_rdy(closest_so_far_out_rsc_rdy_nintersec_loop_one)
    );
  IntersecLoop intersec_loop_two (
      .clk(clk),
      .arst_n(arst_n),
      .quads_rsc_dat(quads_rsc_dat_nintersec_loop_two),
      .quads_rsc_vld(quads_rsc_vld_nintersec_loop_two),
      .quads_rsc_rdy(quads_rsc_rdy_nintersec_loop_two_bud),
      .ray_temp_in_rsc_dat(ray_temp_in_rsc_dat_nintersec_loop_two),
      .ray_temp_in_rsc_vld(ray_temp_in_rsc_vld_nintersec_loop_two),
      .ray_temp_in_rsc_rdy(ray_temp_in_rsc_rdy_nintersec_loop_two_bud),
      .quad_max_in_rsc_dat(quad_max_in_rsc_dat_nintersec_loop_two),
      .quad_max_in_rsc_vld(quad_max_in_rsc_vld_nintersec_loop_two),
      .quad_max_in_rsc_rdy(quad_max_in_rsc_rdy_nintersec_loop_two_bud),
      .quad_hit_anything_out_rsc_dat(quad_hit_anything_out_rsc_dat_nintersec_loop_two),
      .quad_hit_anything_out_rsc_vld(quad_hit_anything_out_rsc_vld_nintersec_loop_two_bud),
      .quad_hit_anything_out_rsc_rdy(quad_hit_anything_out_rsc_rdy_nintersec_loop_two),
      .rec_quad_out_rsc_dat(rec_quad_out_rsc_dat_nintersec_loop_two),
      .rec_quad_out_rsc_vld(rec_quad_out_rsc_vld_nintersec_loop_two_bud),
      .rec_quad_out_rsc_rdy(rec_quad_out_rsc_rdy_nintersec_loop_two),
      .closest_so_far_out_rsc_dat(closest_so_far_out_rsc_dat_nintersec_loop_two),
      .closest_so_far_out_rsc_vld(closest_so_far_out_rsc_vld_nintersec_loop_two_bud),
      .closest_so_far_out_rsc_rdy(closest_so_far_out_rsc_rdy_nintersec_loop_two)
    );
  WorldHit worldHit_1 (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat_nworldHit),
      .ray_in_rsc_vld(ray_in_rsc_vld_nworldHit),
      .ray_in_rsc_rdy(ray_in_rsc_rdy_nworldHit_bud),
      .params_in_rsc_dat(params_in_rsc_dat_nworldHit),
      .params_in_rsc_vld(params_in_rsc_vld_nworldHit),
      .params_in_rsc_rdy(params_in_rsc_rdy_nworldHit_bud),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat_nworldHit),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld_nworldHit),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy_nworldHit_bud),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat_nworldHit),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld_nworldHit),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy_nworldHit_bud),
      .quad_hit_anything_outone_rsc_dat(quad_hit_anything_outone_rsc_dat_nworldHit),
      .quad_hit_anything_outone_rsc_vld(quad_hit_anything_outone_rsc_vld_nworldHit),
      .quad_hit_anything_outone_rsc_rdy(quad_hit_anything_outone_rsc_rdy_nworldHit_bud),
      .quad_hit_anything_outtwo_rsc_dat(quad_hit_anything_outtwo_rsc_dat_nworldHit),
      .quad_hit_anything_outtwo_rsc_vld(quad_hit_anything_outtwo_rsc_vld_nworldHit),
      .quad_hit_anything_outtwo_rsc_rdy(quad_hit_anything_outtwo_rsc_rdy_nworldHit_bud),
      .rec_quad_outone_rsc_dat(rec_quad_outone_rsc_dat_nworldHit),
      .rec_quad_outone_rsc_vld(rec_quad_outone_rsc_vld_nworldHit),
      .rec_quad_outone_rsc_rdy(rec_quad_outone_rsc_rdy_nworldHit_bud),
      .rec_quad_outtwo_rsc_dat(rec_quad_outtwo_rsc_dat_nworldHit),
      .rec_quad_outtwo_rsc_vld(rec_quad_outtwo_rsc_vld_nworldHit),
      .rec_quad_outtwo_rsc_rdy(rec_quad_outtwo_rsc_rdy_nworldHit_bud),
      .closest_so_far_outone_rsc_dat(closest_so_far_outone_rsc_dat_nworldHit),
      .closest_so_far_outone_rsc_vld(closest_so_far_outone_rsc_vld_nworldHit),
      .closest_so_far_outone_rsc_rdy(closest_so_far_outone_rsc_rdy_nworldHit_bud),
      .closest_so_far_outtwo_rsc_dat(closest_so_far_outtwo_rsc_dat_nworldHit),
      .closest_so_far_outtwo_rsc_vld(closest_so_far_outtwo_rsc_vld_nworldHit),
      .closest_so_far_outtwo_rsc_rdy(closest_so_far_outtwo_rsc_rdy_nworldHit_bud),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat_nworldHit),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld_nworldHit_bud),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy_nworldHit),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat_nworldHit),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld_nworldHit_bud),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy_nworldHit),
      .hit_out_rsc_dat(hit_out_rsc_dat_nworldHit),
      .hit_out_rsc_vld(hit_out_rsc_vld_nworldHit_bud),
      .hit_out_rsc_rdy(hit_out_rsc_rdy_nworldHit),
      .ray_out_rsc_dat(ray_out_rsc_dat_nworldHit),
      .ray_out_rsc_vld(ray_out_rsc_vld_nworldHit_bud),
      .ray_out_rsc_rdy(ray_out_rsc_rdy_nworldHit),
      .isHit_rsc_dat(isHit_rsc_dat_nworldHit),
      .isHit_rsc_vld(isHit_rsc_vld_nworldHit_bud),
      .isHit_rsc_rdy(isHit_rsc_rdy_nworldHit)
    );
  MaterialScatter materialScatter_1 (
      .clk(clk),
      .arst_n(arst_n),
      .ray_in_rsc_dat(ray_in_rsc_dat_nmaterialScatter),
      .ray_in_rsc_vld(ray_in_rsc_vld_nmaterialScatter),
      .ray_in_rsc_rdy(ray_in_rsc_rdy_nmaterialScatter_bud),
      .hit_in_rsc_dat(hit_in_rsc_dat_nmaterialScatter),
      .hit_in_rsc_vld(hit_in_rsc_vld_nmaterialScatter),
      .hit_in_rsc_rdy(hit_in_rsc_rdy_nmaterialScatter_bud),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat_nmaterialScatter),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld_nmaterialScatter),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy_nmaterialScatter_bud),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat_nmaterialScatter),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld_nmaterialScatter),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy_nmaterialScatter_bud),
      .isHit_rsc_dat(isHit_rsc_dat_nmaterialScatter),
      .isHit_rsc_vld(isHit_rsc_vld_nmaterialScatter),
      .isHit_rsc_rdy(isHit_rsc_rdy_nmaterialScatter_bud),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat_nmaterialScatter),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld_nmaterialScatter_bud),
      .attenuation_chan_out_rsc_rdy(attenuation_chan_out_rsc_rdy),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat_nmaterialScatter),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld_nmaterialScatter_bud),
      .accumalated_color_out_rsc_rdy(accumalated_color_out_rsc_rdy),
      .ray_out_rsc_dat(ray_out_rsc_dat_nmaterialScatter),
      .ray_out_rsc_vld(ray_out_rsc_vld_nmaterialScatter_bud),
      .ray_out_rsc_rdy(ray_out_rsc_rdy)
    );
  assign ray_in_rsc_rdy = ray_in_rsc_rdy_nloop_distrib_bud;
  assign params_in_rsc_rdy = params_in_rsc_rdy_nloop_distrib_bud;
  assign quad_in_rsc_rdy = quads_rsc_rdy_nloop_distrib_bud;
  assign attenuation_chan_in_rsc_rdy = attenuation_chan_in_rsc_rdy_nloop_distrib_bud;
  assign accumalated_color_chan_in_rsc_rdy = accumalated_color_chan_in_rsc_rdy_nloop_distrib_bud;
  assign attenuation_chan_out_rsc_vld = attenuation_chan_out_rsc_vld_nmaterialScatter_bud;
  assign attenuation_chan_out_rsc_dat = attenuation_chan_out_rsc_dat_nmaterialScatter;
  assign accumalated_color_out_rsc_vld = accumalated_color_out_rsc_vld_nmaterialScatter_bud;
  assign accumalated_color_out_rsc_dat = accumalated_color_out_rsc_dat_nmaterialScatter;
  assign ray_out_rsc_vld = ray_out_rsc_vld_nmaterialScatter_bud;
  assign ray_out_rsc_dat = ray_out_rsc_dat_nmaterialScatter;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ShaderCores
// ------------------------------------------------------------------


module ShaderCores (
  clk, arst_n, quads_in_rsc_dat, quads_in_rsc_vld, quads_in_rsc_rdy, ray_in_rsc_dat,
      ray_in_rsc_vld, ray_in_rsc_rdy, params_in_rsc_dat, params_in_rsc_vld, params_in_rsc_rdy,
      output_pxl_serial_rsc_dat, output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [376:0] quads_in_rsc_dat;
  input quads_in_rsc_vld;
  output quads_in_rsc_rdy;
  input [165:0] ray_in_rsc_dat;
  input ray_in_rsc_vld;
  output ray_in_rsc_rdy;
  input [92:0] params_in_rsc_dat;
  input params_in_rsc_vld;
  output params_in_rsc_rdy;
  output [80:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;


  // Interconnect Declarations
  wire [92:0] params_in_rsc_dat_nshader1;
  wire params_in_rsc_vld_nshader1;
  wire [165:0] ray_in_rsc_dat_nshader1;
  wire ray_in_rsc_vld_nshader1;
  wire [80:0] attenuation_chan_in_rsc_dat_nshader1;
  wire attenuation_chan_in_rsc_vld_nshader1;
  wire [80:0] accumalated_color_chan_in_rsc_dat_nshader1;
  wire accumalated_color_chan_in_rsc_vld_nshader1;
  wire [80:0] attenuation_chan_out_rsc_dat_nshader1;
  wire [80:0] accumalated_color_out_rsc_dat_nshader1;
  wire [165:0] ray_out_rsc_dat_nshader1;
  wire [165:0] ray_scattered_chan_rsc_dat_ncontroller;
  wire ray_scattered_chan_rsc_vld_ncontroller;
  wire [80:0] color_chan_in_rsc_dat_ncontroller;
  wire color_chan_in_rsc_vld_ncontroller;
  wire [80:0] atten_chan_in_rsc_dat_ncontroller;
  wire atten_chan_in_rsc_vld_ncontroller;
  wire [165:0] ray_out_rsc_dat_ncontroller;
  wire ray_out_rsc_rdy_ncontroller;
  wire [92:0] params_out_rsc_dat_ncontroller;
  wire params_out_rsc_rdy_ncontroller;
  wire [80:0] color_chan_out_rsc_dat_ncontroller;
  wire color_chan_out_rsc_rdy_ncontroller;
  wire [80:0] atten_chan_out_rsc_dat_ncontroller;
  wire atten_chan_out_rsc_rdy_ncontroller;
  wire [80:0] output_pxl_serial_rsc_dat_ncontroller;
  wire ray_in_rsc_rdy_nshader1_bud;
  wire ray_out_rsc_vld_ncontroller_bud;
  wire params_in_rsc_rdy_nshader1_bud;
  wire params_out_rsc_vld_ncontroller_bud;
  wire quad_in_rsc_rdy_nshader1_bud;
  wire attenuation_chan_in_rsc_rdy_nshader1_bud;
  wire atten_chan_out_rsc_vld_ncontroller_bud;
  wire accumalated_color_chan_in_rsc_rdy_nshader1_bud;
  wire color_chan_out_rsc_vld_ncontroller_bud;
  wire attenuation_chan_out_rsc_vld_nshader1_bud;
  wire atten_chan_in_rsc_rdy_ncontroller_bud;
  wire accumalated_color_out_rsc_vld_nshader1_bud;
  wire color_chan_in_rsc_rdy_ncontroller_bud;
  wire ray_out_rsc_vld_nshader1_bud;
  wire ray_scattered_chan_rsc_rdy_ncontroller_bud;
  wire ray_chan_in_rsc_rdy_ncontroller_bud;
  wire params_in_rsc_rdy_ncontroller_bud;
  wire output_pxl_serial_rsc_vld_ncontroller_bud;
  wire ray_into_shader_unc_2;
  wire ray_into_shader_idle;
  wire params_to_shader_unc_2;
  wire params_to_shader_idle;
  wire attenuation_chan1_unc_2;
  wire attenuation_chan1_idle;
  wire accumalated_color_chan1_unc_2;
  wire accumalated_color_chan1_idle;
  wire attenuation_chan_out_rsc_rdy_nshader1_prd;
  reg [2:0] attenuation_chan2_cnt;
  wire [3:0] nl_attenuation_chan2_cnt;
  wire attenuation_chan2_prfl;
  wire attenuation_chan2_unc_2;
  wire attenuation_chan2_idle;
  wire accumalated_color_out_rsc_rdy_nshader1_prd;
  reg [2:0] accumalated_color_chan2_cnt;
  wire [3:0] nl_accumalated_color_chan2_cnt;
  wire accumalated_color_chan2_prfl;
  wire accumalated_color_chan2_unc_2;
  wire accumalated_color_chan2_idle;
  wire ray_out_rsc_rdy_nshader1_prd;
  reg [2:0] ray_out1_cnt;
  wire [3:0] nl_ray_out1_cnt;
  wire ray_out1_prfl;
  wire ray_out1_unc_2;
  wire ray_out1_idle;

  wire[0:0] attenuation_chan2_and_3_nl;
  wire[0:0] accumalated_color_chan2_and_3_nl;
  wire[0:0] ray_out1_and_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_attenuation_chan2_cns_pipe_din_vld;
  assign nl_attenuation_chan2_cns_pipe_din_vld = attenuation_chan2_prfl | attenuation_chan_out_rsc_vld_nshader1_bud;
  wire[0:0] attenuation_chan2_not_1_nl;
  wire [80:0] nl_attenuation_chan2_cns_pipe_din;
  assign attenuation_chan2_not_1_nl = ~ attenuation_chan2_prfl;
  assign nl_attenuation_chan2_cns_pipe_din = MUX_v_81_2_2(81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000,
      attenuation_chan_out_rsc_dat_nshader1, (attenuation_chan2_not_1_nl));
  wire [0:0] nl_accumalated_color_chan2_cns_pipe_din_vld;
  assign nl_accumalated_color_chan2_cns_pipe_din_vld = accumalated_color_chan2_prfl
      | accumalated_color_out_rsc_vld_nshader1_bud;
  wire[0:0] accumalated_color_chan2_not_1_nl;
  wire [80:0] nl_accumalated_color_chan2_cns_pipe_din;
  assign accumalated_color_chan2_not_1_nl = ~ accumalated_color_chan2_prfl;
  assign nl_accumalated_color_chan2_cns_pipe_din = MUX_v_81_2_2(81'b000000000000000000000000000000000000000000000000000000000000000000000000000000000,
      accumalated_color_out_rsc_dat_nshader1, (accumalated_color_chan2_not_1_nl));
  wire [0:0] nl_ray_out1_cns_pipe_din_vld;
  assign nl_ray_out1_cns_pipe_din_vld = ray_out1_prfl | ray_out_rsc_vld_nshader1_bud;
  wire[0:0] ray_out1_not_1_nl;
  wire [165:0] nl_ray_out1_cns_pipe_din;
  assign ray_out1_not_1_nl = ~ ray_out1_prfl;
  assign nl_ray_out1_cns_pipe_din = MUX_v_166_2_2(166'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
      ray_out_rsc_dat_nshader1, (ray_out1_not_1_nl));
  wire [0:0] nl_shader1_attenuation_chan_out_rsc_rdy;
  assign nl_shader1_attenuation_chan_out_rsc_rdy = (~ attenuation_chan2_prfl) & attenuation_chan_out_rsc_rdy_nshader1_prd;
  wire [0:0] nl_shader1_accumalated_color_out_rsc_rdy;
  assign nl_shader1_accumalated_color_out_rsc_rdy = (~ accumalated_color_chan2_prfl)
      & accumalated_color_out_rsc_rdy_nshader1_prd;
  wire [0:0] nl_shader1_ray_out_rsc_rdy;
  assign nl_shader1_ray_out_rsc_rdy = (~ ray_out1_prfl) & ray_out_rsc_rdy_nshader1_prd;
  ccs_pipe_v5 #(.rscid(32'sd132),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ray_into_shader_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_rsc_rdy_ncontroller),
      .din_vld(ray_out_rsc_vld_ncontroller_bud),
      .din(ray_out_rsc_dat_ncontroller),
      .dout_rdy(ray_in_rsc_rdy_nshader1_bud),
      .dout_vld(ray_in_rsc_vld_nshader1),
      .dout(ray_in_rsc_dat_nshader1),
      .sz(ray_into_shader_unc_2),
      .sz_req(1'b0),
      .is_idle(ray_into_shader_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd133),
  .width(32'sd93),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) params_to_shader_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(params_out_rsc_rdy_ncontroller),
      .din_vld(params_out_rsc_vld_ncontroller_bud),
      .din(params_out_rsc_dat_ncontroller),
      .dout_rdy(params_in_rsc_rdy_nshader1_bud),
      .dout_vld(params_in_rsc_vld_nshader1),
      .dout(params_in_rsc_dat_nshader1),
      .sz(params_to_shader_unc_2),
      .sz_req(1'b0),
      .is_idle(params_to_shader_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd135),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) attenuation_chan1_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(atten_chan_out_rsc_rdy_ncontroller),
      .din_vld(atten_chan_out_rsc_vld_ncontroller_bud),
      .din(atten_chan_out_rsc_dat_ncontroller),
      .dout_rdy(attenuation_chan_in_rsc_rdy_nshader1_bud),
      .dout_vld(attenuation_chan_in_rsc_vld_nshader1),
      .dout(attenuation_chan_in_rsc_dat_nshader1),
      .sz(attenuation_chan1_unc_2),
      .sz_req(1'b0),
      .is_idle(attenuation_chan1_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd134),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd4),
  .log2_sz(32'sd2),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) accumalated_color_chan1_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(color_chan_out_rsc_rdy_ncontroller),
      .din_vld(color_chan_out_rsc_vld_ncontroller_bud),
      .din(color_chan_out_rsc_dat_ncontroller),
      .dout_rdy(accumalated_color_chan_in_rsc_rdy_nshader1_bud),
      .dout_vld(accumalated_color_chan_in_rsc_vld_nshader1),
      .dout(accumalated_color_chan_in_rsc_dat_nshader1),
      .sz(accumalated_color_chan1_unc_2),
      .sz_req(1'b0),
      .is_idle(accumalated_color_chan1_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd131),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) attenuation_chan2_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(attenuation_chan_out_rsc_rdy_nshader1_prd),
      .din_vld(nl_attenuation_chan2_cns_pipe_din_vld[0:0]),
      .din(nl_attenuation_chan2_cns_pipe_din[80:0]),
      .dout_rdy(atten_chan_in_rsc_rdy_ncontroller_bud),
      .dout_vld(atten_chan_in_rsc_vld_ncontroller),
      .dout(atten_chan_in_rsc_dat_ncontroller),
      .sz(attenuation_chan2_unc_2),
      .sz_req(1'b0),
      .is_idle(attenuation_chan2_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd130),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) accumalated_color_chan2_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(accumalated_color_out_rsc_rdy_nshader1_prd),
      .din_vld(nl_accumalated_color_chan2_cns_pipe_din_vld[0:0]),
      .din(nl_accumalated_color_chan2_cns_pipe_din[80:0]),
      .dout_rdy(color_chan_in_rsc_rdy_ncontroller_bud),
      .dout_vld(color_chan_in_rsc_vld_ncontroller),
      .dout(color_chan_in_rsc_dat_ncontroller),
      .sz(accumalated_color_chan2_unc_2),
      .sz_req(1'b0),
      .is_idle(accumalated_color_chan2_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd129),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ray_out1_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(ray_out_rsc_rdy_nshader1_prd),
      .din_vld(nl_ray_out1_cns_pipe_din_vld[0:0]),
      .din(nl_ray_out1_cns_pipe_din[165:0]),
      .dout_rdy(ray_scattered_chan_rsc_rdy_ncontroller_bud),
      .dout_vld(ray_scattered_chan_rsc_vld_ncontroller),
      .dout(ray_scattered_chan_rsc_dat_ncontroller),
      .sz(ray_out1_unc_2),
      .sz_req(1'b0),
      .is_idle(ray_out1_idle)
    );
  Shader shader1 (
      .clk(clk),
      .arst_n(arst_n),
      .params_in_rsc_dat(params_in_rsc_dat_nshader1),
      .params_in_rsc_vld(params_in_rsc_vld_nshader1),
      .params_in_rsc_rdy(params_in_rsc_rdy_nshader1_bud),
      .quad_in_rsc_dat(quads_in_rsc_dat),
      .quad_in_rsc_vld(quads_in_rsc_vld),
      .quad_in_rsc_rdy(quad_in_rsc_rdy_nshader1_bud),
      .ray_in_rsc_dat(ray_in_rsc_dat_nshader1),
      .ray_in_rsc_vld(ray_in_rsc_vld_nshader1),
      .ray_in_rsc_rdy(ray_in_rsc_rdy_nshader1_bud),
      .attenuation_chan_in_rsc_dat(attenuation_chan_in_rsc_dat_nshader1),
      .attenuation_chan_in_rsc_vld(attenuation_chan_in_rsc_vld_nshader1),
      .attenuation_chan_in_rsc_rdy(attenuation_chan_in_rsc_rdy_nshader1_bud),
      .accumalated_color_chan_in_rsc_dat(accumalated_color_chan_in_rsc_dat_nshader1),
      .accumalated_color_chan_in_rsc_vld(accumalated_color_chan_in_rsc_vld_nshader1),
      .accumalated_color_chan_in_rsc_rdy(accumalated_color_chan_in_rsc_rdy_nshader1_bud),
      .attenuation_chan_out_rsc_dat(attenuation_chan_out_rsc_dat_nshader1),
      .attenuation_chan_out_rsc_vld(attenuation_chan_out_rsc_vld_nshader1_bud),
      .attenuation_chan_out_rsc_rdy(nl_shader1_attenuation_chan_out_rsc_rdy[0:0]),
      .accumalated_color_out_rsc_dat(accumalated_color_out_rsc_dat_nshader1),
      .accumalated_color_out_rsc_vld(accumalated_color_out_rsc_vld_nshader1_bud),
      .accumalated_color_out_rsc_rdy(nl_shader1_accumalated_color_out_rsc_rdy[0:0]),
      .ray_out_rsc_dat(ray_out_rsc_dat_nshader1),
      .ray_out_rsc_vld(ray_out_rsc_vld_nshader1_bud),
      .ray_out_rsc_rdy(nl_shader1_ray_out_rsc_rdy[0:0])
    );
  ShaderFeedbackController controller (
      .clk(clk),
      .arst_n(arst_n),
      .ray_chan_in_rsc_dat(ray_in_rsc_dat),
      .ray_chan_in_rsc_vld(ray_in_rsc_vld),
      .ray_chan_in_rsc_rdy(ray_chan_in_rsc_rdy_ncontroller_bud),
      .ray_scattered_chan_rsc_dat(ray_scattered_chan_rsc_dat_ncontroller),
      .ray_scattered_chan_rsc_vld(ray_scattered_chan_rsc_vld_ncontroller),
      .ray_scattered_chan_rsc_rdy(ray_scattered_chan_rsc_rdy_ncontroller_bud),
      .params_in_rsc_dat(params_in_rsc_dat),
      .params_in_rsc_vld(params_in_rsc_vld),
      .params_in_rsc_rdy(params_in_rsc_rdy_ncontroller_bud),
      .color_chan_in_rsc_dat(color_chan_in_rsc_dat_ncontroller),
      .color_chan_in_rsc_vld(color_chan_in_rsc_vld_ncontroller),
      .color_chan_in_rsc_rdy(color_chan_in_rsc_rdy_ncontroller_bud),
      .atten_chan_in_rsc_dat(atten_chan_in_rsc_dat_ncontroller),
      .atten_chan_in_rsc_vld(atten_chan_in_rsc_vld_ncontroller),
      .atten_chan_in_rsc_rdy(atten_chan_in_rsc_rdy_ncontroller_bud),
      .ray_out_rsc_dat(ray_out_rsc_dat_ncontroller),
      .ray_out_rsc_vld(ray_out_rsc_vld_ncontroller_bud),
      .ray_out_rsc_rdy(ray_out_rsc_rdy_ncontroller),
      .params_out_rsc_dat(params_out_rsc_dat_ncontroller),
      .params_out_rsc_vld(params_out_rsc_vld_ncontroller_bud),
      .params_out_rsc_rdy(params_out_rsc_rdy_ncontroller),
      .color_chan_out_rsc_dat(color_chan_out_rsc_dat_ncontroller),
      .color_chan_out_rsc_vld(color_chan_out_rsc_vld_ncontroller_bud),
      .color_chan_out_rsc_rdy(color_chan_out_rsc_rdy_ncontroller),
      .atten_chan_out_rsc_dat(atten_chan_out_rsc_dat_ncontroller),
      .atten_chan_out_rsc_vld(atten_chan_out_rsc_vld_ncontroller_bud),
      .atten_chan_out_rsc_rdy(atten_chan_out_rsc_rdy_ncontroller),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat_ncontroller),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld_ncontroller_bud),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy)
    );
  assign quads_in_rsc_rdy = quad_in_rsc_rdy_nshader1_bud;
  assign attenuation_chan2_prfl = ~((attenuation_chan2_cnt==3'b100));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      attenuation_chan2_cnt <= 3'b000;
    end
    else begin
      attenuation_chan2_cnt <= nl_attenuation_chan2_cnt[2:0];
    end
  end
  assign attenuation_chan2_and_3_nl = attenuation_chan2_prfl & attenuation_chan_out_rsc_rdy_nshader1_prd;
  assign nl_attenuation_chan2_cnt  = attenuation_chan2_cnt + conv_u2u_1_3(attenuation_chan2_and_3_nl);
  assign accumalated_color_chan2_prfl = ~((accumalated_color_chan2_cnt==3'b100));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      accumalated_color_chan2_cnt <= 3'b000;
    end
    else begin
      accumalated_color_chan2_cnt <= nl_accumalated_color_chan2_cnt[2:0];
    end
  end
  assign accumalated_color_chan2_and_3_nl = accumalated_color_chan2_prfl & accumalated_color_out_rsc_rdy_nshader1_prd;
  assign nl_accumalated_color_chan2_cnt  = accumalated_color_chan2_cnt + conv_u2u_1_3(accumalated_color_chan2_and_3_nl);
  assign ray_out1_prfl = ~((ray_out1_cnt==3'b100));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ray_out1_cnt <= 3'b000;
    end
    else begin
      ray_out1_cnt <= nl_ray_out1_cnt[2:0];
    end
  end
  assign ray_out1_and_3_nl = ray_out1_prfl & ray_out_rsc_rdy_nshader1_prd;
  assign nl_ray_out1_cnt  = ray_out1_cnt + conv_u2u_1_3(ray_out1_and_3_nl);
  assign ray_in_rsc_rdy = ray_chan_in_rsc_rdy_ncontroller_bud;
  assign params_in_rsc_rdy = params_in_rsc_rdy_ncontroller_bud;
  assign output_pxl_serial_rsc_vld = output_pxl_serial_rsc_vld_ncontroller_bud;
  assign output_pxl_serial_rsc_dat = output_pxl_serial_rsc_dat_ncontroller;

  function automatic [165:0] MUX_v_166_2_2;
    input [165:0] input_0;
    input [165:0] input_1;
    input [0:0] sel;
    reg [165:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_166_2_2 = result;
  end
  endfunction


  function automatic [80:0] MUX_v_81_2_2;
    input [80:0] input_0;
    input [80:0] input_1;
    input [0:0] sel;
    reg [80:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_81_2_2 = result;
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    RendererWrapper
// ------------------------------------------------------------------


module RendererWrapper (
  clk, arst_n, quads_in_rsc_dat, quads_in_rsc_vld, quads_in_rsc_rdy, render_params_rsc_dat,
      render_params_rsc_vld, render_params_rsc_rdy, output_pxl_sample_rsc_dat, output_pxl_sample_rsc_vld,
      output_pxl_sample_rsc_rdy
);
  input clk;
  input arst_n;
  input [376:0] quads_in_rsc_dat;
  input quads_in_rsc_vld;
  output quads_in_rsc_rdy;
  input [419:0] render_params_rsc_dat;
  input render_params_rsc_vld;
  output render_params_rsc_rdy;
  output [80:0] output_pxl_sample_rsc_dat;
  output output_pxl_sample_rsc_vld;
  input output_pxl_sample_rsc_rdy;


  // Interconnect Declarations
  wire [419:0] render_params_out_rsc_dat_nrenderLooper;
  wire render_params_out_rsc_rdy_nrenderLooper;
  wire [22:0] loopIndicesOut_rsc_dat_nrenderLooper;
  wire loopIndicesOut_rsc_rdy_nrenderLooper;
  wire [22:0] loopIndicesIn_rsc_dat_nrayGeneration;
  wire loopIndicesIn_rsc_vld_nrayGeneration;
  wire [419:0] paramsIn_rsc_dat_nrayGeneration;
  wire paramsIn_rsc_vld_nrayGeneration;
  wire [92:0] paramsOut_rsc_dat_nrayGeneration;
  wire paramsOut_rsc_rdy_nrayGeneration;
  wire [165:0] rayOut_rsc_dat_nrayGeneration;
  wire rayOut_rsc_rdy_nrayGeneration;
  wire [165:0] ray_in_rsc_dat_nshaderCores;
  wire ray_in_rsc_vld_nshaderCores;
  wire [92:0] params_in_rsc_dat_nshaderCores;
  wire params_in_rsc_vld_nshaderCores;
  wire [80:0] output_pxl_serial_rsc_dat_nshaderCores;
  wire [165:0] rayIn_rsc_dat_nrayCollector;
  wire rayIn_rsc_vld_nrayCollector;
  wire [92:0] paramsIn_rsc_dat_nrayCollector;
  wire paramsIn_rsc_vld_nrayCollector;
  wire [92:0] paramsOut_rsc_dat_nrayCollector;
  wire paramsOut_rsc_rdy_nrayCollector;
  wire [165:0] rayOut_rsc_dat_nrayCollector;
  wire rayOut_rsc_rdy_nrayCollector;
  wire render_params_rsc_rdy_nrenderLooper_bud;
  wire render_params_out_rsc_vld_nrenderLooper_bud;
  wire paramsIn_rsc_rdy_nrayGeneration_bud;
  wire loopIndicesOut_rsc_vld_nrenderLooper_bud;
  wire loopIndicesIn_rsc_rdy_nrayGeneration_bud;
  wire paramsOut_rsc_vld_nrayGeneration_bud;
  wire paramsIn_rsc_rdy_nrayCollector_bud;
  wire rayOut_rsc_vld_nrayGeneration_bud;
  wire rayIn_rsc_rdy_nrayCollector_bud;
  wire quads_in_rsc_rdy_nshaderCores_bud;
  wire ray_in_rsc_rdy_nshaderCores_bud;
  wire rayOut_rsc_vld_nrayCollector_bud;
  wire params_in_rsc_rdy_nshaderCores_bud;
  wire paramsOut_rsc_vld_nrayCollector_bud;
  wire output_pxl_serial_rsc_vld_nshaderCores_bud;
  wire paramsChanneltoRayGen_unc_2;
  wire paramsChanneltoRayGen_idle;
  wire loopIndicesChanneltoRayGen_unc_2;
  wire loopIndicesChanneltoRayGen_idle;
  wire paramsChanneltoCollector_unc_2;
  wire paramsChanneltoCollector_idle;
  wire rayOut_unc_2;
  wire rayOut_idle;
  wire rayToShader_unc_2;
  wire rayToShader_idle;
  wire paramsChanneltoShader_unc_2;
  wire paramsChanneltoShader_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd145),
  .width(32'sd420),
  .sz_width(32'sd1),
  .fifo_sz(32'sd5),
  .log2_sz(32'sd3),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) paramsChanneltoRayGen_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(render_params_out_rsc_rdy_nrenderLooper),
      .din_vld(render_params_out_rsc_vld_nrenderLooper_bud),
      .din(render_params_out_rsc_dat_nrenderLooper),
      .dout_rdy(paramsIn_rsc_rdy_nrayGeneration_bud),
      .dout_vld(paramsIn_rsc_vld_nrayGeneration),
      .dout(paramsIn_rsc_dat_nrayGeneration),
      .sz(paramsChanneltoRayGen_unc_2),
      .sz_req(1'b0),
      .is_idle(paramsChanneltoRayGen_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd148),
  .width(32'sd23),
  .sz_width(32'sd1),
  .fifo_sz(32'sd5),
  .log2_sz(32'sd3),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) loopIndicesChanneltoRayGen_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(loopIndicesOut_rsc_rdy_nrenderLooper),
      .din_vld(loopIndicesOut_rsc_vld_nrenderLooper_bud),
      .din(loopIndicesOut_rsc_dat_nrenderLooper),
      .dout_rdy(loopIndicesIn_rsc_rdy_nrayGeneration_bud),
      .dout_vld(loopIndicesIn_rsc_vld_nrayGeneration),
      .dout(loopIndicesIn_rsc_dat_nrayGeneration),
      .sz(loopIndicesChanneltoRayGen_unc_2),
      .sz_req(1'b0),
      .is_idle(loopIndicesChanneltoRayGen_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd146),
  .width(32'sd93),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) paramsChanneltoCollector_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(paramsOut_rsc_rdy_nrayGeneration),
      .din_vld(paramsOut_rsc_vld_nrayGeneration_bud),
      .din(paramsOut_rsc_dat_nrayGeneration),
      .dout_rdy(paramsIn_rsc_rdy_nrayCollector_bud),
      .dout_vld(paramsIn_rsc_vld_nrayCollector),
      .dout(paramsIn_rsc_dat_nrayCollector),
      .sz(paramsChanneltoCollector_unc_2),
      .sz_req(1'b0),
      .is_idle(paramsChanneltoCollector_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd143),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayOut_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(rayOut_rsc_rdy_nrayGeneration),
      .din_vld(rayOut_rsc_vld_nrayGeneration_bud),
      .din(rayOut_rsc_dat_nrayGeneration),
      .dout_rdy(rayIn_rsc_rdy_nrayCollector_bud),
      .dout_vld(rayIn_rsc_vld_nrayCollector),
      .dout(rayIn_rsc_dat_nrayCollector),
      .sz(rayOut_unc_2),
      .sz_req(1'b0),
      .is_idle(rayOut_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd144),
  .width(32'sd166),
  .sz_width(32'sd1),
  .fifo_sz(32'sd18),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) rayToShader_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(rayOut_rsc_rdy_nrayCollector),
      .din_vld(rayOut_rsc_vld_nrayCollector_bud),
      .din(rayOut_rsc_dat_nrayCollector),
      .dout_rdy(ray_in_rsc_rdy_nshaderCores_bud),
      .dout_vld(ray_in_rsc_vld_nshaderCores),
      .dout(ray_in_rsc_dat_nshaderCores),
      .sz(rayToShader_unc_2),
      .sz_req(1'b0),
      .is_idle(rayToShader_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd147),
  .width(32'sd93),
  .sz_width(32'sd1),
  .fifo_sz(32'sd18),
  .log2_sz(32'sd5),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) paramsChanneltoShader_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(paramsOut_rsc_rdy_nrayCollector),
      .din_vld(paramsOut_rsc_vld_nrayCollector_bud),
      .din(paramsOut_rsc_dat_nrayCollector),
      .dout_rdy(params_in_rsc_rdy_nshaderCores_bud),
      .dout_vld(params_in_rsc_vld_nshaderCores),
      .dout(params_in_rsc_dat_nshaderCores),
      .sz(paramsChanneltoShader_unc_2),
      .sz_req(1'b0),
      .is_idle(paramsChanneltoShader_idle)
    );
  RenderLooper renderLooper_1 (
      .clk(clk),
      .arst_n(arst_n),
      .render_params_rsc_dat(render_params_rsc_dat),
      .render_params_rsc_vld(render_params_rsc_vld),
      .render_params_rsc_rdy(render_params_rsc_rdy_nrenderLooper_bud),
      .render_params_out_rsc_dat(render_params_out_rsc_dat_nrenderLooper),
      .render_params_out_rsc_vld(render_params_out_rsc_vld_nrenderLooper_bud),
      .render_params_out_rsc_rdy(render_params_out_rsc_rdy_nrenderLooper),
      .loopIndicesOut_rsc_dat(loopIndicesOut_rsc_dat_nrenderLooper),
      .loopIndicesOut_rsc_vld(loopIndicesOut_rsc_vld_nrenderLooper_bud),
      .loopIndicesOut_rsc_rdy(loopIndicesOut_rsc_rdy_nrenderLooper)
    );
  RayGeneration rayGeneration_1 (
      .clk(clk),
      .arst_n(arst_n),
      .loopIndicesIn_rsc_dat(loopIndicesIn_rsc_dat_nrayGeneration),
      .loopIndicesIn_rsc_vld(loopIndicesIn_rsc_vld_nrayGeneration),
      .loopIndicesIn_rsc_rdy(loopIndicesIn_rsc_rdy_nrayGeneration_bud),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nrayGeneration),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nrayGeneration),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nrayGeneration_bud),
      .paramsOut_rsc_dat(paramsOut_rsc_dat_nrayGeneration),
      .paramsOut_rsc_vld(paramsOut_rsc_vld_nrayGeneration_bud),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy_nrayGeneration),
      .rayOut_rsc_dat(rayOut_rsc_dat_nrayGeneration),
      .rayOut_rsc_vld(rayOut_rsc_vld_nrayGeneration_bud),
      .rayOut_rsc_rdy(rayOut_rsc_rdy_nrayGeneration)
    );
  ShaderCores shaderCores_1 (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsc_dat(quads_in_rsc_dat),
      .quads_in_rsc_vld(quads_in_rsc_vld),
      .quads_in_rsc_rdy(quads_in_rsc_rdy_nshaderCores_bud),
      .ray_in_rsc_dat(ray_in_rsc_dat_nshaderCores),
      .ray_in_rsc_vld(ray_in_rsc_vld_nshaderCores),
      .ray_in_rsc_rdy(ray_in_rsc_rdy_nshaderCores_bud),
      .params_in_rsc_dat(params_in_rsc_dat_nshaderCores),
      .params_in_rsc_vld(params_in_rsc_vld_nshaderCores),
      .params_in_rsc_rdy(params_in_rsc_rdy_nshaderCores_bud),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat_nshaderCores),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld_nshaderCores_bud),
      .output_pxl_serial_rsc_rdy(output_pxl_sample_rsc_rdy)
    );
  RayCollector rayCollector_1 (
      .clk(clk),
      .arst_n(arst_n),
      .rayIn_rsc_dat(rayIn_rsc_dat_nrayCollector),
      .rayIn_rsc_vld(rayIn_rsc_vld_nrayCollector),
      .rayIn_rsc_rdy(rayIn_rsc_rdy_nrayCollector_bud),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nrayCollector),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nrayCollector),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nrayCollector_bud),
      .paramsOut_rsc_dat(paramsOut_rsc_dat_nrayCollector),
      .paramsOut_rsc_vld(paramsOut_rsc_vld_nrayCollector_bud),
      .paramsOut_rsc_rdy(paramsOut_rsc_rdy_nrayCollector),
      .rayOut_rsc_dat(rayOut_rsc_dat_nrayCollector),
      .rayOut_rsc_vld(rayOut_rsc_vld_nrayCollector_bud),
      .rayOut_rsc_rdy(rayOut_rsc_rdy_nrayCollector)
    );
  assign render_params_rsc_rdy = render_params_rsc_rdy_nrenderLooper_bud;
  assign quads_in_rsc_rdy = quads_in_rsc_rdy_nshaderCores_bud;
  assign output_pxl_sample_rsc_vld = output_pxl_serial_rsc_vld_nshaderCores_bud;
  assign output_pxl_sample_rsc_dat = output_pxl_serial_rsc_dat_nshaderCores;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Pathtracer_struct
// ------------------------------------------------------------------


module Pathtracer_struct (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      output_pxl_serial_rsc_dat_b, output_pxl_serial_rsc_dat_g, output_pxl_serial_rsc_dat_r,
      output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [11:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [7:0] output_pxl_serial_rsc_dat_b;
  output [7:0] output_pxl_serial_rsc_dat_g;
  output [7:0] output_pxl_serial_rsc_dat_r;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;


  // Interconnect Declarations
  wire [56:0] qbuffer_params_rsc_dat_nparamsDeserializer;
  wire qbuffer_params_rsc_rdy_nparamsDeserializer;
  wire [419:0] render_params_rsc_dat_nparamsDeserializer;
  wire render_params_rsc_rdy_nparamsDeserializer;
  wire [419:0] accum_params_rsc_dat_nparamsDeserializer;
  wire accum_params_rsc_rdy_nparamsDeserializer;
  wire [376:0] quad_serial_out_rsc_dat_nparamsDeserializer;
  wire quad_serial_out_rsc_rdy_nparamsDeserializer;
  wire [376:0] quads_in_rsc_dat_nquadsBuffer;
  wire quads_in_rsc_vld_nquadsBuffer;
  wire [56:0] paramsIn_rsc_dat_nquadsBuffer;
  wire paramsIn_rsc_vld_nquadsBuffer;
  wire [376:0] quads_out_rsc_dat_nquadsBuffer;
  wire quads_out_rsc_rdy_nquadsBuffer;
  wire [376:0] quads_in_rsc_dat_nrenderer;
  wire quads_in_rsc_vld_nrenderer;
  wire [419:0] render_params_rsc_dat_nrenderer;
  wire render_params_rsc_vld_nrenderer;
  wire [80:0] output_pxl_sample_rsc_dat_nrenderer;
  wire output_pxl_sample_rsc_rdy_nrenderer;
  wire [419:0] accumulator_parms_rsc_dat_npixelAccumulator;
  wire accumulator_parms_rsc_vld_npixelAccumulator;
  wire [80:0] pxl_sample_rsc_dat_npixelAccumulator;
  wire pxl_sample_rsc_vld_npixelAccumulator;
  wire [23:0] output_pxl_serial_rsc_dat_npixelAccumulator;
  wire inputChannel_rsc_rdy_nparamsDeserializer_bud;
  wire qbuffer_params_rsc_vld_nparamsDeserializer_bud;
  wire paramsIn_rsc_rdy_nquadsBuffer_bud;
  wire render_params_rsc_vld_nparamsDeserializer_bud;
  wire render_params_rsc_rdy_nrenderer_bud;
  wire accum_params_rsc_vld_nparamsDeserializer_bud;
  wire accumulator_parms_rsc_rdy_npixelAccumulator_bud;
  wire quad_serial_out_rsc_vld_nparamsDeserializer_bud;
  wire quads_in_rsc_rdy_nquadsBuffer_bud;
  wire quads_out_rsc_vld_nquadsBuffer_bud;
  wire quads_in_rsc_rdy_nrenderer_bud;
  wire output_pxl_sample_rsc_vld_nrenderer_bud;
  wire pxl_sample_rsc_rdy_npixelAccumulator_bud;
  wire output_pxl_serial_rsc_vld_npixelAccumulator_bud;
  wire quad_buffer_params_unc_2;
  wire quad_buffer_params_idle;
  wire renderer_params_unc_2;
  wire renderer_params_idle;
  wire accumulator_params_unc_2;
  wire accumulator_params_idle;
  wire quad_serial_unc_2;
  wire quad_serial_idle;
  wire quads_out_unc_2;
  wire quads_out_idle;
  wire pxl_sample_unc_2;
  wire pxl_sample_idle;


  // Interconnect Declarations for Component Instantiations 
  ccs_pipe_v5 #(.rscid(32'sd158),
  .width(32'sd57),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_buffer_params_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(qbuffer_params_rsc_rdy_nparamsDeserializer),
      .din_vld(qbuffer_params_rsc_vld_nparamsDeserializer_bud),
      .din(qbuffer_params_rsc_dat_nparamsDeserializer),
      .dout_rdy(paramsIn_rsc_rdy_nquadsBuffer_bud),
      .dout_vld(paramsIn_rsc_vld_nquadsBuffer),
      .dout(paramsIn_rsc_dat_nquadsBuffer),
      .sz(quad_buffer_params_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_buffer_params_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd156),
  .width(32'sd420),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) renderer_params_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(render_params_rsc_rdy_nparamsDeserializer),
      .din_vld(render_params_rsc_vld_nparamsDeserializer_bud),
      .din(render_params_rsc_dat_nparamsDeserializer),
      .dout_rdy(render_params_rsc_rdy_nrenderer_bud),
      .dout_vld(render_params_rsc_vld_nrenderer),
      .dout(render_params_rsc_dat_nrenderer),
      .sz(renderer_params_unc_2),
      .sz_req(1'b0),
      .is_idle(renderer_params_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd157),
  .width(32'sd420),
  .sz_width(32'sd1),
  .fifo_sz(32'sd1),
  .log2_sz(32'sd0),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) accumulator_params_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(accum_params_rsc_rdy_nparamsDeserializer),
      .din_vld(accum_params_rsc_vld_nparamsDeserializer_bud),
      .din(accum_params_rsc_dat_nparamsDeserializer),
      .dout_rdy(accumulator_parms_rsc_rdy_npixelAccumulator_bud),
      .dout_vld(accumulator_parms_rsc_vld_npixelAccumulator),
      .dout(accumulator_parms_rsc_dat_npixelAccumulator),
      .sz(accumulator_params_unc_2),
      .sz_req(1'b0),
      .is_idle(accumulator_params_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd154),
  .width(32'sd377),
  .sz_width(32'sd1),
  .fifo_sz(32'sd125),
  .log2_sz(32'sd7),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quad_serial_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quad_serial_out_rsc_rdy_nparamsDeserializer),
      .din_vld(quad_serial_out_rsc_vld_nparamsDeserializer_bud),
      .din(quad_serial_out_rsc_dat_nparamsDeserializer),
      .dout_rdy(quads_in_rsc_rdy_nquadsBuffer_bud),
      .dout_vld(quads_in_rsc_vld_nquadsBuffer),
      .dout(quads_in_rsc_dat_nquadsBuffer),
      .sz(quad_serial_unc_2),
      .sz_req(1'b0),
      .is_idle(quad_serial_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd155),
  .width(32'sd377),
  .sz_width(32'sd1),
  .fifo_sz(32'sd7),
  .log2_sz(32'sd3),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) quads_out_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(quads_out_rsc_rdy_nquadsBuffer),
      .din_vld(quads_out_rsc_vld_nquadsBuffer_bud),
      .din(quads_out_rsc_dat_nquadsBuffer),
      .dout_rdy(quads_in_rsc_rdy_nrenderer_bud),
      .dout_vld(quads_in_rsc_vld_nrenderer),
      .dout(quads_in_rsc_dat_nrenderer),
      .sz(quads_out_unc_2),
      .sz_req(1'b0),
      .is_idle(quads_out_idle)
    );
  ccs_pipe_v5 #(.rscid(32'sd159),
  .width(32'sd81),
  .sz_width(32'sd1),
  .fifo_sz(32'sd2),
  .log2_sz(32'sd1),
  .ph_clk(32'sd1),
  .ph_en(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) pxl_sample_cns_pipe (
      .clk(clk),
      .en(1'b0),
      .arst(arst_n),
      .srst(1'b1),
      .din_rdy(output_pxl_sample_rsc_rdy_nrenderer),
      .din_vld(output_pxl_sample_rsc_vld_nrenderer_bud),
      .din(output_pxl_sample_rsc_dat_nrenderer),
      .dout_rdy(pxl_sample_rsc_rdy_npixelAccumulator_bud),
      .dout_vld(pxl_sample_rsc_vld_npixelAccumulator),
      .dout(pxl_sample_rsc_dat_npixelAccumulator),
      .sz(pxl_sample_unc_2),
      .sz_req(1'b0),
      .is_idle(pxl_sample_idle)
    );
  ParamsDeserializer paramsDeserializer_1 (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy_nparamsDeserializer_bud),
      .qbuffer_params_rsc_dat(qbuffer_params_rsc_dat_nparamsDeserializer),
      .qbuffer_params_rsc_vld(qbuffer_params_rsc_vld_nparamsDeserializer_bud),
      .qbuffer_params_rsc_rdy(qbuffer_params_rsc_rdy_nparamsDeserializer),
      .render_params_rsc_dat(render_params_rsc_dat_nparamsDeserializer),
      .render_params_rsc_vld(render_params_rsc_vld_nparamsDeserializer_bud),
      .render_params_rsc_rdy(render_params_rsc_rdy_nparamsDeserializer),
      .accum_params_rsc_dat(accum_params_rsc_dat_nparamsDeserializer),
      .accum_params_rsc_vld(accum_params_rsc_vld_nparamsDeserializer_bud),
      .accum_params_rsc_rdy(accum_params_rsc_rdy_nparamsDeserializer),
      .quad_serial_out_rsc_dat(quad_serial_out_rsc_dat_nparamsDeserializer),
      .quad_serial_out_rsc_vld(quad_serial_out_rsc_vld_nparamsDeserializer_bud),
      .quad_serial_out_rsc_rdy(quad_serial_out_rsc_rdy_nparamsDeserializer)
    );
  QuadBuffer_64 quadsBuffer (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsc_dat(quads_in_rsc_dat_nquadsBuffer),
      .quads_in_rsc_vld(quads_in_rsc_vld_nquadsBuffer),
      .quads_in_rsc_rdy(quads_in_rsc_rdy_nquadsBuffer_bud),
      .paramsIn_rsc_dat(paramsIn_rsc_dat_nquadsBuffer),
      .paramsIn_rsc_vld(paramsIn_rsc_vld_nquadsBuffer),
      .paramsIn_rsc_rdy(paramsIn_rsc_rdy_nquadsBuffer_bud),
      .quads_out_rsc_dat(quads_out_rsc_dat_nquadsBuffer),
      .quads_out_rsc_vld(quads_out_rsc_vld_nquadsBuffer_bud),
      .quads_out_rsc_rdy(quads_out_rsc_rdy_nquadsBuffer)
    );
  RendererWrapper renderer (
      .clk(clk),
      .arst_n(arst_n),
      .quads_in_rsc_dat(quads_in_rsc_dat_nrenderer),
      .quads_in_rsc_vld(quads_in_rsc_vld_nrenderer),
      .quads_in_rsc_rdy(quads_in_rsc_rdy_nrenderer_bud),
      .render_params_rsc_dat(render_params_rsc_dat_nrenderer),
      .render_params_rsc_vld(render_params_rsc_vld_nrenderer),
      .render_params_rsc_rdy(render_params_rsc_rdy_nrenderer_bud),
      .output_pxl_sample_rsc_dat(output_pxl_sample_rsc_dat_nrenderer),
      .output_pxl_sample_rsc_vld(output_pxl_sample_rsc_vld_nrenderer_bud),
      .output_pxl_sample_rsc_rdy(output_pxl_sample_rsc_rdy_nrenderer)
    );
  PixelAccumulator pixelAccumulator_1 (
      .clk(clk),
      .arst_n(arst_n),
      .accumulator_parms_rsc_dat(accumulator_parms_rsc_dat_npixelAccumulator),
      .accumulator_parms_rsc_vld(accumulator_parms_rsc_vld_npixelAccumulator),
      .accumulator_parms_rsc_rdy(accumulator_parms_rsc_rdy_npixelAccumulator_bud),
      .pxl_sample_rsc_dat(pxl_sample_rsc_dat_npixelAccumulator),
      .pxl_sample_rsc_vld(pxl_sample_rsc_vld_npixelAccumulator),
      .pxl_sample_rsc_rdy(pxl_sample_rsc_rdy_npixelAccumulator_bud),
      .output_pxl_serial_rsc_dat(output_pxl_serial_rsc_dat_npixelAccumulator),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld_npixelAccumulator_bud),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy)
    );
  assign output_pxl_serial_rsc_dat_r = output_pxl_serial_rsc_dat_npixelAccumulator[7:0];
  assign output_pxl_serial_rsc_dat_g = output_pxl_serial_rsc_dat_npixelAccumulator[15:8];
  assign output_pxl_serial_rsc_dat_b = output_pxl_serial_rsc_dat_npixelAccumulator[23:16];
  assign inputChannel_rsc_rdy = inputChannel_rsc_rdy_nparamsDeserializer_bud;
  assign output_pxl_serial_rsc_vld = output_pxl_serial_rsc_vld_npixelAccumulator_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Pathtracer
// ------------------------------------------------------------------


module Pathtracer (
  clk, arst_n, inputChannel_rsc_dat, inputChannel_rsc_vld, inputChannel_rsc_rdy,
      output_pxl_serial_rsc_dat, output_pxl_serial_rsc_vld, output_pxl_serial_rsc_rdy
);
  input clk;
  input arst_n;
  input [11:0] inputChannel_rsc_dat;
  input inputChannel_rsc_vld;
  output inputChannel_rsc_rdy;
  output [23:0] output_pxl_serial_rsc_dat;
  output output_pxl_serial_rsc_vld;
  input output_pxl_serial_rsc_rdy;


  // Interconnect Declarations
  wire [7:0] output_pxl_serial_rsc_dat_b;
  wire [7:0] output_pxl_serial_rsc_dat_g;
  wire [7:0] output_pxl_serial_rsc_dat_r;


  // Interconnect Declarations for Component Instantiations 
  Pathtracer_struct Pathtracer_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .inputChannel_rsc_dat(inputChannel_rsc_dat),
      .inputChannel_rsc_vld(inputChannel_rsc_vld),
      .inputChannel_rsc_rdy(inputChannel_rsc_rdy),
      .output_pxl_serial_rsc_dat_b(output_pxl_serial_rsc_dat_b),
      .output_pxl_serial_rsc_dat_g(output_pxl_serial_rsc_dat_g),
      .output_pxl_serial_rsc_dat_r(output_pxl_serial_rsc_dat_r),
      .output_pxl_serial_rsc_vld(output_pxl_serial_rsc_vld),
      .output_pxl_serial_rsc_rdy(output_pxl_serial_rsc_rdy)
    );
  assign output_pxl_serial_rsc_dat = {output_pxl_serial_rsc_dat_b , output_pxl_serial_rsc_dat_g
      , output_pxl_serial_rsc_dat_r};
endmodule



